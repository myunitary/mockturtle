// Benchmark "/tmp/tmp" written by ABC on Sat Nov  8 22:34:36 2025

module Lite_MIPS_firstframe ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128, po129, po130, po131, po132, po133, po134, po135, po136,
    po137, po138, po139, po140, po141, po142, po143, po144, po145, po146,
    po147, po148, po149, po150, po151, po152, po153, po154, po155, po156,
    po157, po158, po159, po160, po161, po162, po163, po164, po165, po166,
    po167, po168, po169, po170, po171, po172, po173, po174, po175, po176,
    po177, po178, po179, po180, po181, po182, po183, po184, po185, po186,
    po187, po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215, po216,
    po217, po218, po219, po220, po221, po222, po223, po224, po225, po226,
    po227, po228, po229, po230, po231, po232, po233, po234, po235, po236,
    po237, po238, po239, po240, po241, po242, po243, po244, po245, po246,
    po247, po248, po249, po250, po251, po252, po253, po254, po255, po256,
    po257, po258, po259, po260, po261, po262, po263, po264, po265, po266,
    po267, po268, po269, po270, po271, po272, po273, po274, po275, po276,
    po277, po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305, po306,
    po307, po308, po309, po310, po311, po312, po313, po314, po315, po316,
    po317, po318, po319, po320, po321, po322, po323, po324, po325, po326,
    po327, po328, po329, po330, po331, po332, po333, po334, po335, po336,
    po337, po338, po339, po340, po341, po342, po343, po344, po345, po346,
    po347, po348, po349, po350, po351, po352, po353, po354, po355, po356,
    po357, po358, po359, po360, po361, po362, po363, po364, po365, po366,
    po367, po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395, po396,
    po397, po398, po399, po400, po401, po402, po403, po404, po405, po406,
    po407, po408, po409, po410, po411, po412, po413, po414, po415, po416,
    po417, po418, po419, po420, po421, po422, po423, po424, po425, po426,
    po427, po428, po429, po430, po431, po432, po433, po434, po435, po436,
    po437, po438, po439, po440, po441, po442, po443, po444, po445, po446,
    po447, po448, po449, po450, po451, po452, po453, po454, po455, po456,
    po457, po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485, po486,
    po487, po488, po489, po490, po491, po492, po493, po494, po495, po496,
    po497, po498, po499, po500, po501, po502, po503, po504, po505, po506,
    po507, po508, po509, po510, po511, po512, po513, po514, po515, po516,
    po517, po518, po519, po520, po521, po522, po523, po524, po525, po526,
    po527, po528, po529, po530, po531, po532, po533, po534, po535, po536,
    po537, po538, po539, po540, po541, po542, po543, po544, po545, po546,
    po547, po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575, po576,
    po577, po578, po579, po580, po581, po582, po583, po584, po585, po586,
    po587, po588, po589, po590, po591, po592, po593, po594, po595, po596,
    po597, po598, po599, po600, po601, po602, po603, po604, po605, po606,
    po607, po608, po609, po610, po611, po612, po613, po614, po615, po616,
    po617, po618, po619, po620, po621, po622, po623, po624, po625, po626,
    po627, po628, po629, po630, po631, po632, po633, po634, po635, po636,
    po637, po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665, po666,
    po667, po668, po669, po670, po671, po672, po673, po674, po675, po676,
    po677, po678, po679, po680, po681, po682, po683, po684, po685, po686,
    po687, po688, po689, po690, po691, po692, po693, po694, po695, po696,
    po697, po698, po699, po700, po701, po702, po703, po704, po705, po706,
    po707, po708, po709, po710, po711, po712, po713, po714, po715, po716,
    po717, po718, po719, po720, po721, po722, po723, po724, po725, po726,
    po727, po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755, po756,
    po757, po758, po759, po760, po761, po762, po763, po764, po765, po766,
    po767, po768, po769, po770, po771, po772, po773, po774, po775, po776,
    po777, po778, po779, po780, po781, po782, po783, po784, po785, po786,
    po787, po788, po789, po790, po791, po792, po793, po794, po795, po796,
    po797, po798, po799, po800, po801, po802, po803, po804, po805, po806,
    po807, po808, po809, po810, po811, po812, po813, po814, po815, po816,
    po817, po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845, po846,
    po847, po848, po849, po850, po851, po852, po853, po854, po855, po856,
    po857, po858, po859, po860, po861, po862, po863, po864, po865, po866,
    po867, po868, po869, po870, po871, po872, po873, po874, po875, po876,
    po877, po878, po879, po880, po881, po882, po883, po884, po885, po886,
    po887, po888, po889, po890, po891, po892, po893, po894, po895, po896,
    po897, po898, po899, po900, po901, po902, po903, po904, po905, po906,
    po907, po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935, po936,
    po937, po938, po939, po940, po941, po942, po943, po944, po945, po946,
    po947, po948, po949, po950, po951, po952, po953, po954, po955, po956,
    po957, po958, po959, po960, po961, po962, po963, po964, po965, po966,
    po967, po968, po969, po970, po971, po972, po973, po974, po975, po976,
    po977, po978, po979, po980, po981, po982, po983, po984, po985, po986,
    po987, po988, po989, po990, po991, po992, po993, po994, po995, po996,
    po997, po998, po999, po1000, po1001, po1002, po1003, po1004, po1005,
    po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014,
    po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023,
    po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032,
    po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041,
    po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050,
    po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059,
    po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068,
    po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077,
    po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086,
    po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095,
    po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104,
    po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113,
    po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122,
    po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131,
    po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140,
    po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149,
    po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158,
    po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167,
    po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176,
    po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185,
    po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194,
    po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203,
    po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212,
    po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221,
    po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230,
    po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239,
    po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248,
    po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257,
    po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266,
    po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275,
    po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284,
    po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293,
    po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302,
    po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311,
    po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320,
    po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329,
    po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338,
    po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347,
    po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356,
    po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365,
    po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374,
    po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383,
    po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392,
    po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401,
    po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410,
    po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419,
    po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428,
    po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437,
    po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446,
    po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455,
    po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464,
    po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473,
    po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482,
    po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491,
    po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500,
    po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509,
    po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518,
    po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527,
    po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536,
    po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545,
    po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554,
    po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563,
    po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572,
    po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581,
    po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590,
    po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599,
    po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608,
    po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617,
    po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626,
    po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635,
    po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644,
    po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653,
    po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662,
    po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671,
    po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680,
    po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689,
    po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698,
    po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707,
    po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716,
    po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725,
    po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734,
    po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743,
    po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752,
    po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761,
    po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770,
    po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779,
    po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788,
    po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797,
    po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806,
    po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815,
    po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824,
    po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833,
    po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842,
    po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851,
    po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860,
    po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869,
    po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878,
    po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887,
    po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896,
    po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905,
    po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914,
    po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923,
    po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932,
    po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941,
    po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950,
    po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959,
    po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968,
    po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977,
    po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986,
    po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995,
    po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004,
    po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013,
    po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022,
    po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031,
    po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040,
    po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049,
    po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058,
    po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067,
    po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076,
    po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085,
    po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094,
    po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103,
    po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112,
    po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121,
    po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130,
    po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139,
    po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148,
    po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157,
    po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166,
    po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175,
    po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184,
    po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193,
    po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202,
    po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211,
    po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220,
    po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229,
    po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238,
    po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247,
    po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256,
    po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265,
    po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274,
    po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283,
    po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292,
    po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301,
    po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310,
    po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319,
    po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328,
    po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337,
    po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346,
    po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355,
    po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364,
    po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373,
    po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382,
    po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391,
    po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400,
    po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409,
    po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418,
    po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427,
    po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436,
    po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445,
    po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454,
    po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463,
    po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472,
    po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481,
    po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490,
    po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499,
    po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508,
    po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517,
    po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526,
    po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535,
    po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544,
    po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553,
    po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562,
    po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571,
    po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580,
    po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589,
    po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598,
    po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607,
    po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616,
    po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625,
    po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634,
    po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643,
    po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652,
    po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661,
    po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670,
    po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679,
    po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688,
    po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697,
    po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706,
    po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715,
    po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724,
    po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733,
    po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742,
    po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751,
    po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760,
    po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769,
    po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778,
    po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787,
    po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796,
    po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805,
    po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814,
    po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823,
    po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832,
    po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841,
    po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850,
    po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859,
    po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868,
    po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877,
    po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886,
    po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895,
    po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904,
    po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913,
    po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922,
    po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931,
    po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940,
    po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949,
    po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958,
    po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967,
    po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976,
    po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985,
    po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994,
    po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003,
    po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012,
    po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021,
    po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030,
    po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039,
    po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048,
    po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057,
    po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066,
    po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075,
    po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084,
    po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093,
    po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102,
    po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111,
    po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120,
    po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129,
    po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138,
    po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147,
    po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156,
    po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165,
    po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174,
    po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183,
    po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192,
    po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201,
    po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210,
    po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219,
    po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228,
    po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237,
    po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246,
    po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255,
    po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264,
    po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273,
    po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282,
    po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291,
    po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300,
    po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309,
    po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318,
    po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327,
    po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336,
    po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345,
    po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354,
    po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363,
    po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372,
    po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381,
    po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390,
    po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399,
    po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408,
    po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417,
    po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426,
    po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435,
    po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444,
    po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453,
    po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462,
    po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471,
    po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480,
    po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489,
    po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498,
    po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507,
    po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516,
    po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525,
    po3526, po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534,
    po3535, po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543,
    po3544, po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552,
    po3553, po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561,
    po3562, po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570,
    po3571, po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579,
    po3580, po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588,
    po3589, po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597,
    po3598, po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606,
    po3607, po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615,
    po3616, po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624,
    po3625, po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633,
    po3634, po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642,
    po3643, po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651,
    po3652, po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660,
    po3661, po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669,
    po3670, po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678,
    po3679, po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687,
    po3688, po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696,
    po3697, po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705,
    po3706, po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714,
    po3715, po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723,
    po3724, po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732,
    po3733, po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741,
    po3742, po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750,
    po3751, po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759,
    po3760, po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768,
    po3769, po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777,
    po3778, po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786,
    po3787, po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795,
    po3796, po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804,
    po3805, po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813,
    po3814, po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822,
    po3823, po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831,
    po3832, po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840,
    po3841, po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849,
    po3850, po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858,
    po3859, po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867,
    po3868, po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876,
    po3877, po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885,
    po3886, po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894,
    po3895, po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903,
    po3904, po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912,
    po3913, po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921,
    po3922, po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930,
    po3931, po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939,
    po3940, po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948,
    po3949, po3950, po3951, po3952, po3953, po3954, po3955, po3956, po3957,
    po3958, po3959, po3960, po3961, po3962, po3963, po3964, po3965, po3966,
    po3967, po3968, po3969, po3970, po3971, po3972, po3973, po3974, po3975,
    po3976, po3977, po3978, po3979, po3980, po3981, po3982, po3983, po3984,
    po3985, po3986, po3987, po3988, po3989, po3990, po3991, po3992, po3993,
    po3994, po3995, po3996, po3997, po3998, po3999, po4000, po4001, po4002,
    po4003, po4004, po4005, po4006, po4007, po4008, po4009, po4010, po4011,
    po4012, po4013, po4014, po4015, po4016, po4017, po4018, po4019, po4020,
    po4021, po4022, po4023, po4024, po4025, po4026, po4027, po4028, po4029,
    po4030, po4031, po4032, po4033, po4034, po4035, po4036, po4037, po4038,
    po4039, po4040, po4041, po4042, po4043, po4044, po4045, po4046, po4047,
    po4048, po4049, po4050, po4051, po4052, po4053, po4054, po4055, po4056,
    po4057, po4058, po4059, po4060, po4061, po4062, po4063, po4064, po4065,
    po4066, po4067, po4068, po4069, po4070, po4071, po4072, po4073, po4074,
    po4075, po4076, po4077, po4078, po4079, po4080, po4081, po4082, po4083,
    po4084, po4085, po4086, po4087, po4088, po4089, po4090, po4091, po4092,
    po4093, po4094, po4095, po4096, po4097, po4098, po4099, po4100, po4101,
    po4102, po4103, po4104, po4105, po4106, po4107, po4108, po4109, po4110,
    po4111, po4112, po4113, po4114, po4115, po4116, po4117, po4118, po4119,
    po4120, po4121, po4122, po4123, po4124, po4125, po4126, po4127, po4128,
    po4129, po4130, po4131, po4132, po4133, po4134, po4135, po4136, po4137,
    po4138, po4139, po4140, po4141, po4142, po4143, po4144, po4145, po4146,
    po4147, po4148, po4149, po4150, po4151, po4152, po4153, po4154, po4155,
    po4156, po4157, po4158, po4159, po4160, po4161, po4162, po4163, po4164,
    po4165, po4166, po4167, po4168, po4169, po4170, po4171, po4172, po4173,
    po4174, po4175, po4176, po4177, po4178, po4179, po4180, po4181, po4182,
    po4183, po4184, po4185, po4186, po4187, po4188, po4189, po4190, po4191,
    po4192, po4193, po4194, po4195, po4196, po4197, po4198, po4199, po4200,
    po4201, po4202, po4203, po4204, po4205, po4206, po4207, po4208, po4209,
    po4210, po4211, po4212, po4213, po4214, po4215, po4216, po4217, po4218,
    po4219, po4220, po4221, po4222, po4223, po4224, po4225, po4226, po4227,
    po4228, po4229, po4230, po4231, po4232, po4233, po4234, po4235, po4236,
    po4237, po4238, po4239, po4240, po4241, po4242, po4243, po4244, po4245,
    po4246, po4247, po4248, po4249, po4250, po4251, po4252, po4253, po4254,
    po4255, po4256, po4257, po4258, po4259, po4260, po4261, po4262, po4263,
    po4264, po4265, po4266, po4267, po4268, po4269, po4270, po4271, po4272,
    po4273, po4274, po4275, po4276, po4277, po4278, po4279, po4280, po4281,
    po4282, po4283, po4284, po4285, po4286, po4287, po4288, po4289, po4290,
    po4291, po4292, po4293, po4294, po4295, po4296, po4297, po4298, po4299,
    po4300, po4301, po4302, po4303, po4304, po4305, po4306, po4307, po4308,
    po4309, po4310, po4311, po4312, po4313, po4314, po4315, po4316, po4317,
    po4318, po4319, po4320, po4321, po4322, po4323, po4324, po4325, po4326,
    po4327, po4328, po4329, po4330, po4331, po4332, po4333, po4334, po4335,
    po4336, po4337, po4338, po4339, po4340, po4341, po4342, po4343, po4344,
    po4345, po4346, po4347, po4348, po4349, po4350, po4351, po4352, po4353,
    po4354, po4355, po4356, po4357, po4358, po4359, po4360, po4361, po4362,
    po4363, po4364, po4365, po4366, po4367, po4368, po4369, po4370, po4371,
    po4372, po4373, po4374, po4375, po4376, po4377, po4378, po4379, po4380,
    po4381, po4382, po4383, po4384, po4385, po4386, po4387, po4388, po4389,
    po4390, po4391, po4392, po4393, po4394, po4395, po4396, po4397, po4398,
    po4399, po4400, po4401, po4402, po4403, po4404, po4405, po4406, po4407,
    po4408, po4409, po4410, po4411, po4412, po4413, po4414, po4415, po4416,
    po4417, po4418, po4419, po4420, po4421, po4422, po4423, po4424, po4425,
    po4426, po4427, po4428, po4429, po4430, po4431, po4432, po4433, po4434,
    po4435, po4436, po4437, po4438, po4439, po4440, po4441, po4442, po4443,
    po4444, po4445, po4446, po4447, po4448, po4449, po4450, po4451, po4452,
    po4453, po4454, po4455, po4456, po4457, po4458, po4459, po4460, po4461,
    po4462, po4463, po4464, po4465, po4466, po4467, po4468, po4469, po4470,
    po4471, po4472, po4473, po4474, po4475, po4476, po4477, po4478, po4479,
    po4480, po4481, po4482, po4483, po4484, po4485, po4486, po4487, po4488,
    po4489, po4490, po4491, po4492, po4493, po4494, po4495, po4496, po4497,
    po4498, po4499, po4500, po4501, po4502, po4503, po4504, po4505, po4506,
    po4507, po4508, po4509, po4510, po4511, po4512, po4513, po4514, po4515,
    po4516, po4517, po4518, po4519, po4520, po4521, po4522, po4523, po4524,
    po4525, po4526, po4527, po4528, po4529, po4530, po4531, po4532, po4533,
    po4534, po4535, po4536, po4537, po4538, po4539, po4540, po4541, po4542,
    po4543, po4544, po4545, po4546, po4547, po4548, po4549, po4550, po4551,
    po4552, po4553, po4554, po4555, po4556, po4557, po4558, po4559, po4560,
    po4561, po4562, po4563, po4564, po4565, po4566, po4567, po4568, po4569,
    po4570, po4571, po4572, po4573, po4574, po4575, po4576, po4577, po4578,
    po4579, po4580, po4581, po4582, po4583, po4584, po4585, po4586, po4587,
    po4588, po4589, po4590, po4591, po4592, po4593, po4594, po4595, po4596,
    po4597, po4598, po4599, po4600, po4601, po4602, po4603, po4604, po4605,
    po4606, po4607, po4608, po4609, po4610, po4611, po4612, po4613, po4614,
    po4615, po4616, po4617, po4618, po4619, po4620, po4621, po4622, po4623,
    po4624, po4625, po4626, po4627, po4628, po4629, po4630, po4631, po4632,
    po4633, po4634, po4635, po4636, po4637, po4638, po4639, po4640, po4641,
    po4642, po4643, po4644, po4645, po4646, po4647, po4648, po4649, po4650,
    po4651, po4652, po4653, po4654, po4655, po4656, po4657, po4658, po4659,
    po4660, po4661, po4662, po4663, po4664, po4665, po4666, po4667, po4668,
    po4669, po4670, po4671, po4672, po4673, po4674, po4675, po4676, po4677,
    po4678, po4679, po4680, po4681, po4682, po4683, po4684, po4685, po4686,
    po4687, po4688, po4689, po4690, po4691, po4692, po4693, po4694, po4695,
    po4696, po4697, po4698, po4699, po4700, po4701, po4702, po4703, po4704,
    po4705, po4706, po4707, po4708, po4709, po4710, po4711, po4712, po4713,
    po4714, po4715, po4716, po4717, po4718, po4719, po4720, po4721, po4722,
    po4723, po4724, po4725, po4726, po4727, po4728, po4729, po4730, po4731,
    po4732, po4733, po4734, po4735, po4736, po4737, po4738, po4739, po4740,
    po4741, po4742, po4743, po4744, po4745, po4746, po4747, po4748, po4749,
    po4750, po4751, po4752, po4753, po4754, po4755, po4756, po4757, po4758,
    po4759, po4760, po4761, po4762, po4763, po4764, po4765, po4766, po4767,
    po4768, po4769, po4770, po4771, po4772, po4773, po4774, po4775, po4776,
    po4777, po4778, po4779, po4780, po4781, po4782, po4783, po4784, po4785,
    po4786, po4787, po4788, po4789, po4790, po4791, po4792, po4793, po4794,
    po4795, po4796, po4797, po4798, po4799, po4800, po4801, po4802, po4803,
    po4804, po4805, po4806, po4807, po4808, po4809, po4810, po4811, po4812,
    po4813, po4814, po4815, po4816, po4817, po4818, po4819, po4820, po4821,
    po4822, po4823, po4824, po4825, po4826, po4827, po4828, po4829, po4830,
    po4831, po4832, po4833, po4834, po4835, po4836, po4837, po4838, po4839,
    po4840, po4841, po4842, po4843, po4844, po4845, po4846, po4847, po4848,
    po4849, po4850, po4851, po4852, po4853, po4854, po4855, po4856, po4857,
    po4858, po4859, po4860, po4861, po4862, po4863, po4864, po4865, po4866,
    po4867, po4868, po4869, po4870, po4871, po4872, po4873, po4874, po4875,
    po4876, po4877, po4878, po4879, po4880, po4881, po4882, po4883, po4884,
    po4885, po4886, po4887, po4888, po4889, po4890, po4891, po4892, po4893,
    po4894, po4895, po4896, po4897, po4898, po4899, po4900, po4901, po4902,
    po4903, po4904, po4905, po4906, po4907, po4908, po4909, po4910, po4911,
    po4912, po4913, po4914, po4915, po4916, po4917, po4918, po4919, po4920,
    po4921, po4922, po4923, po4924, po4925, po4926, po4927, po4928, po4929,
    po4930, po4931, po4932, po4933, po4934, po4935, po4936, po4937, po4938,
    po4939, po4940, po4941, po4942, po4943, po4944, po4945, po4946, po4947,
    po4948, po4949, po4950, po4951, po4952, po4953, po4954, po4955, po4956,
    po4957, po4958, po4959, po4960, po4961, po4962, po4963, po4964, po4965,
    po4966, po4967, po4968, po4969, po4970, po4971, po4972, po4973, po4974,
    po4975, po4976, po4977, po4978, po4979, po4980, po4981, po4982, po4983,
    po4984, po4985, po4986, po4987, po4988, po4989, po4990, po4991, po4992,
    po4993, po4994, po4995, po4996, po4997, po4998, po4999, po5000, po5001,
    po5002, po5003, po5004, po5005, po5006, po5007, po5008, po5009, po5010,
    po5011, po5012, po5013, po5014, po5015, po5016, po5017, po5018, po5019,
    po5020, po5021, po5022, po5023, po5024, po5025, po5026, po5027, po5028,
    po5029, po5030, po5031, po5032, po5033, po5034, po5035, po5036, po5037,
    po5038, po5039, po5040, po5041, po5042, po5043, po5044, po5045, po5046,
    po5047, po5048, po5049, po5050, po5051, po5052, po5053, po5054, po5055,
    po5056, po5057, po5058, po5059, po5060, po5061, po5062, po5063, po5064,
    po5065, po5066, po5067, po5068, po5069, po5070, po5071, po5072, po5073,
    po5074, po5075, po5076, po5077, po5078, po5079, po5080, po5081, po5082,
    po5083, po5084, po5085, po5086, po5087, po5088, po5089, po5090, po5091,
    po5092, po5093, po5094, po5095, po5096, po5097, po5098, po5099, po5100,
    po5101, po5102, po5103, po5104, po5105, po5106, po5107, po5108, po5109,
    po5110, po5111, po5112, po5113, po5114, po5115, po5116, po5117, po5118,
    po5119, po5120, po5121, po5122, po5123, po5124, po5125, po5126, po5127,
    po5128, po5129, po5130, po5131, po5132, po5133, po5134, po5135, po5136,
    po5137, po5138, po5139, po5140, po5141, po5142, po5143, po5144, po5145,
    po5146, po5147, po5148, po5149, po5150, po5151, po5152, po5153, po5154,
    po5155, po5156, po5157, po5158, po5159, po5160, po5161, po5162, po5163,
    po5164, po5165, po5166, po5167, po5168, po5169, po5170, po5171, po5172,
    po5173, po5174, po5175, po5176, po5177, po5178, po5179, po5180, po5181,
    po5182, po5183, po5184, po5185, po5186, po5187, po5188, po5189, po5190,
    po5191, po5192, po5193, po5194, po5195, po5196, po5197, po5198, po5199,
    po5200, po5201, po5202, po5203, po5204, po5205, po5206, po5207, po5208,
    po5209, po5210, po5211, po5212, po5213, po5214, po5215, po5216, po5217,
    po5218, po5219, po5220, po5221, po5222, po5223, po5224, po5225, po5226,
    po5227, po5228, po5229, po5230, po5231, po5232, po5233, po5234, po5235,
    po5236, po5237, po5238, po5239, po5240, po5241, po5242, po5243, po5244,
    po5245, po5246, po5247, po5248, po5249, po5250, po5251, po5252, po5253,
    po5254, po5255, po5256, po5257, po5258, po5259, po5260, po5261, po5262,
    po5263, po5264, po5265, po5266, po5267, po5268, po5269, po5270, po5271,
    po5272, po5273, po5274, po5275, po5276, po5277, po5278, po5279, po5280,
    po5281, po5282, po5283, po5284, po5285, po5286, po5287, po5288, po5289,
    po5290, po5291, po5292, po5293, po5294, po5295, po5296, po5297, po5298,
    po5299, po5300, po5301, po5302, po5303, po5304, po5305, po5306, po5307,
    po5308, po5309, po5310, po5311, po5312, po5313, po5314, po5315, po5316,
    po5317, po5318, po5319, po5320, po5321, po5322, po5323, po5324, po5325,
    po5326, po5327, po5328, po5329, po5330, po5331, po5332, po5333, po5334,
    po5335, po5336, po5337, po5338, po5339, po5340, po5341, po5342, po5343,
    po5344, po5345, po5346, po5347, po5348, po5349, po5350, po5351, po5352,
    po5353, po5354, po5355, po5356, po5357, po5358, po5359, po5360, po5361,
    po5362, po5363, po5364, po5365, po5366, po5367, po5368, po5369, po5370,
    po5371, po5372, po5373, po5374, po5375, po5376, po5377, po5378, po5379,
    po5380, po5381, po5382, po5383, po5384, po5385, po5386, po5387, po5388,
    po5389, po5390, po5391, po5392, po5393, po5394, po5395, po5396, po5397,
    po5398, po5399, po5400, po5401, po5402, po5403, po5404, po5405, po5406,
    po5407, po5408, po5409, po5410, po5411, po5412, po5413, po5414, po5415,
    po5416, po5417, po5418, po5419, po5420, po5421, po5422, po5423, po5424,
    po5425, po5426, po5427, po5428, po5429, po5430, po5431, po5432, po5433,
    po5434, po5435, po5436, po5437, po5438, po5439, po5440, po5441, po5442,
    po5443, po5444, po5445, po5446, po5447, po5448, po5449, po5450, po5451,
    po5452, po5453, po5454, po5455, po5456, po5457, po5458, po5459, po5460,
    po5461, po5462, po5463, po5464, po5465, po5466, po5467, po5468, po5469,
    po5470, po5471, po5472, po5473, po5474, po5475, po5476, po5477, po5478,
    po5479, po5480, po5481, po5482, po5483, po5484, po5485, po5486, po5487,
    po5488, po5489, po5490, po5491, po5492, po5493, po5494, po5495, po5496,
    po5497, po5498, po5499, po5500, po5501, po5502, po5503, po5504, po5505,
    po5506, po5507, po5508, po5509, po5510, po5511, po5512, po5513, po5514,
    po5515, po5516, po5517, po5518, po5519, po5520, po5521, po5522, po5523,
    po5524, po5525, po5526, po5527, po5528, po5529, po5530, po5531, po5532,
    po5533, po5534, po5535, po5536, po5537, po5538, po5539, po5540, po5541,
    po5542, po5543, po5544, po5545, po5546, po5547, po5548, po5549, po5550,
    po5551, po5552, po5553, po5554, po5555, po5556, po5557, po5558, po5559,
    po5560, po5561, po5562, po5563, po5564, po5565, po5566, po5567, po5568,
    po5569, po5570, po5571, po5572, po5573, po5574, po5575, po5576, po5577,
    po5578, po5579, po5580, po5581, po5582, po5583, po5584, po5585, po5586,
    po5587, po5588, po5589, po5590, po5591, po5592, po5593, po5594, po5595,
    po5596, po5597, po5598, po5599, po5600, po5601, po5602, po5603, po5604,
    po5605, po5606, po5607, po5608, po5609, po5610, po5611, po5612, po5613,
    po5614, po5615, po5616, po5617, po5618, po5619, po5620, po5621, po5622,
    po5623, po5624, po5625, po5626, po5627, po5628, po5629, po5630, po5631,
    po5632, po5633, po5634, po5635, po5636, po5637, po5638, po5639, po5640,
    po5641, po5642, po5643, po5644, po5645, po5646, po5647, po5648, po5649,
    po5650, po5651, po5652, po5653, po5654, po5655, po5656, po5657, po5658,
    po5659, po5660, po5661, po5662, po5663, po5664, po5665, po5666, po5667,
    po5668, po5669, po5670, po5671, po5672, po5673, po5674, po5675, po5676,
    po5677, po5678, po5679, po5680, po5681, po5682, po5683, po5684, po5685,
    po5686, po5687, po5688, po5689, po5690, po5691, po5692, po5693, po5694,
    po5695, po5696, po5697, po5698, po5699, po5700, po5701, po5702, po5703,
    po5704, po5705, po5706, po5707, po5708, po5709, po5710, po5711, po5712,
    po5713, po5714, po5715, po5716, po5717, po5718, po5719, po5720, po5721,
    po5722, po5723, po5724, po5725, po5726, po5727, po5728, po5729, po5730,
    po5731, po5732, po5733, po5734, po5735, po5736, po5737, po5738, po5739,
    po5740, po5741, po5742, po5743, po5744, po5745, po5746, po5747, po5748,
    po5749, po5750, po5751, po5752, po5753, po5754, po5755, po5756, po5757,
    po5758, po5759, po5760, po5761, po5762, po5763, po5764, po5765, po5766,
    po5767, po5768, po5769, po5770, po5771, po5772, po5773, po5774, po5775,
    po5776, po5777, po5778, po5779, po5780, po5781, po5782, po5783, po5784,
    po5785, po5786, po5787, po5788, po5789, po5790, po5791, po5792, po5793,
    po5794, po5795, po5796, po5797, po5798, po5799, po5800, po5801, po5802,
    po5803, po5804, po5805, po5806, po5807, po5808, po5809, po5810, po5811,
    po5812, po5813, po5814, po5815, po5816, po5817, po5818, po5819, po5820,
    po5821, po5822, po5823, po5824, po5825, po5826, po5827, po5828, po5829,
    po5830, po5831, po5832, po5833, po5834, po5835, po5836, po5837, po5838,
    po5839, po5840, po5841, po5842, po5843, po5844, po5845, po5846, po5847,
    po5848, po5849, po5850, po5851, po5852, po5853, po5854, po5855, po5856,
    po5857, po5858, po5859, po5860, po5861, po5862, po5863, po5864, po5865,
    po5866, po5867, po5868, po5869, po5870, po5871, po5872, po5873, po5874,
    po5875, po5876, po5877, po5878, po5879, po5880, po5881, po5882, po5883,
    po5884, po5885, po5886, po5887, po5888, po5889, po5890, po5891, po5892,
    po5893, po5894, po5895, po5896, po5897, po5898, po5899, po5900, po5901,
    po5902, po5903, po5904, po5905, po5906, po5907, po5908, po5909, po5910,
    po5911, po5912, po5913, po5914, po5915, po5916, po5917, po5918, po5919,
    po5920, po5921, po5922, po5923, po5924, po5925, po5926, po5927, po5928,
    po5929, po5930, po5931, po5932, po5933, po5934, po5935, po5936, po5937,
    po5938, po5939, po5940, po5941, po5942, po5943, po5944, po5945, po5946,
    po5947, po5948, po5949, po5950, po5951, po5952, po5953, po5954, po5955,
    po5956, po5957, po5958, po5959, po5960, po5961, po5962, po5963, po5964,
    po5965, po5966, po5967, po5968, po5969, po5970, po5971, po5972, po5973,
    po5974, po5975, po5976, po5977, po5978, po5979, po5980, po5981, po5982,
    po5983, po5984, po5985, po5986, po5987, po5988, po5989, po5990, po5991,
    po5992, po5993, po5994, po5995, po5996, po5997, po5998, po5999, po6000,
    po6001, po6002, po6003, po6004, po6005, po6006, po6007, po6008, po6009,
    po6010, po6011, po6012, po6013, po6014, po6015, po6016, po6017, po6018,
    po6019, po6020, po6021, po6022, po6023, po6024, po6025, po6026, po6027,
    po6028, po6029, po6030, po6031, po6032, po6033, po6034, po6035, po6036,
    po6037, po6038, po6039, po6040, po6041, po6042, po6043, po6044, po6045,
    po6046, po6047, po6048, po6049, po6050, po6051, po6052, po6053, po6054,
    po6055, po6056, po6057, po6058, po6059, po6060, po6061, po6062, po6063,
    po6064, po6065, po6066, po6067, po6068, po6069, po6070, po6071, po6072,
    po6073, po6074, po6075, po6076, po6077, po6078, po6079, po6080, po6081,
    po6082, po6083, po6084, po6085, po6086, po6087, po6088, po6089, po6090,
    po6091, po6092, po6093, po6094, po6095, po6096, po6097, po6098, po6099,
    po6100, po6101, po6102, po6103, po6104, po6105, po6106, po6107, po6108,
    po6109, po6110, po6111, po6112, po6113, po6114, po6115, po6116, po6117,
    po6118, po6119, po6120, po6121, po6122, po6123, po6124, po6125, po6126,
    po6127, po6128, po6129, po6130, po6131, po6132, po6133, po6134, po6135,
    po6136, po6137, po6138, po6139, po6140, po6141, po6142, po6143, po6144,
    po6145, po6146, po6147, po6148, po6149, po6150, po6151, po6152, po6153,
    po6154, po6155, po6156, po6157, po6158, po6159, po6160, po6161, po6162,
    po6163, po6164, po6165, po6166, po6167, po6168, po6169, po6170, po6171,
    po6172, po6173, po6174, po6175, po6176, po6177, po6178, po6179, po6180,
    po6181, po6182, po6183, po6184, po6185, po6186, po6187, po6188, po6189,
    po6190, po6191, po6192, po6193, po6194, po6195, po6196, po6197, po6198,
    po6199, po6200, po6201, po6202, po6203, po6204, po6205, po6206, po6207,
    po6208, po6209, po6210, po6211, po6212, po6213, po6214, po6215, po6216,
    po6217, po6218, po6219, po6220, po6221, po6222, po6223, po6224, po6225,
    po6226, po6227, po6228, po6229, po6230, po6231, po6232, po6233, po6234,
    po6235, po6236, po6237, po6238, po6239, po6240, po6241, po6242, po6243,
    po6244, po6245, po6246, po6247, po6248, po6249, po6250, po6251, po6252,
    po6253, po6254, po6255, po6256, po6257, po6258, po6259, po6260, po6261,
    po6262, po6263, po6264, po6265, po6266, po6267, po6268, po6269, po6270,
    po6271, po6272, po6273, po6274, po6275, po6276, po6277, po6278, po6279,
    po6280, po6281, po6282, po6283, po6284, po6285, po6286, po6287, po6288,
    po6289, po6290, po6291, po6292, po6293, po6294, po6295, po6296, po6297,
    po6298, po6299, po6300, po6301, po6302, po6303, po6304, po6305, po6306,
    po6307, po6308, po6309, po6310, po6311, po6312, po6313, po6314, po6315,
    po6316, po6317, po6318, po6319, po6320, po6321, po6322, po6323, po6324,
    po6325, po6326, po6327, po6328, po6329, po6330, po6331, po6332, po6333,
    po6334, po6335, po6336, po6337, po6338, po6339, po6340, po6341, po6342,
    po6343, po6344, po6345, po6346, po6347, po6348, po6349, po6350, po6351,
    po6352, po6353, po6354, po6355, po6356, po6357, po6358, po6359, po6360,
    po6361, po6362, po6363, po6364, po6365, po6366, po6367, po6368, po6369,
    po6370, po6371, po6372, po6373, po6374, po6375, po6376, po6377, po6378,
    po6379, po6380, po6381, po6382, po6383, po6384, po6385, po6386, po6387,
    po6388, po6389, po6390, po6391, po6392, po6393, po6394, po6395, po6396,
    po6397, po6398, po6399, po6400, po6401, po6402, po6403, po6404, po6405,
    po6406, po6407, po6408, po6409, po6410, po6411, po6412, po6413, po6414,
    po6415, po6416, po6417, po6418, po6419, po6420, po6421, po6422, po6423,
    po6424, po6425, po6426, po6427, po6428, po6429, po6430, po6431, po6432,
    po6433, po6434, po6435, po6436, po6437, po6438, po6439, po6440, po6441,
    po6442, po6443, po6444, po6445, po6446, po6447, po6448, po6449, po6450,
    po6451, po6452, po6453, po6454, po6455, po6456, po6457, po6458, po6459,
    po6460, po6461, po6462, po6463, po6464, po6465, po6466, po6467, po6468,
    po6469, po6470, po6471, po6472, po6473, po6474, po6475, po6476, po6477,
    po6478, po6479, po6480, po6481, po6482, po6483, po6484, po6485, po6486,
    po6487, po6488, po6489, po6490, po6491, po6492, po6493, po6494, po6495,
    po6496, po6497, po6498, po6499, po6500, po6501, po6502, po6503, po6504,
    po6505, po6506, po6507, po6508, po6509, po6510, po6511, po6512, po6513,
    po6514, po6515, po6516, po6517, po6518, po6519, po6520, po6521, po6522,
    po6523, po6524, po6525, po6526, po6527, po6528, po6529, po6530, po6531,
    po6532, po6533, po6534, po6535, po6536, po6537, po6538, po6539, po6540,
    po6541, po6542, po6543, po6544, po6545, po6546, po6547, po6548, po6549,
    po6550, po6551, po6552, po6553, po6554, po6555, po6556, po6557, po6558,
    po6559, po6560, po6561, po6562, po6563, po6564, po6565, po6566, po6567,
    po6568, po6569, po6570, po6571, po6572, po6573, po6574, po6575, po6576,
    po6577, po6578, po6579, po6580, po6581, po6582, po6583, po6584, po6585,
    po6586, po6587, po6588, po6589, po6590, po6591, po6592, po6593, po6594,
    po6595, po6596, po6597, po6598, po6599, po6600, po6601, po6602, po6603,
    po6604, po6605, po6606, po6607, po6608, po6609, po6610, po6611, po6612,
    po6613, po6614, po6615, po6616, po6617, po6618, po6619, po6620, po6621,
    po6622, po6623, po6624, po6625, po6626, po6627, po6628, po6629, po6630,
    po6631, po6632, po6633, po6634, po6635, po6636, po6637, po6638, po6639,
    po6640, po6641, po6642, po6643, po6644, po6645, po6646, po6647, po6648,
    po6649, po6650, po6651, po6652, po6653, po6654, po6655, po6656, po6657,
    po6658, po6659, po6660, po6661, po6662, po6663, po6664, po6665, po6666,
    po6667, po6668, po6669, po6670, po6671, po6672, po6673, po6674, po6675,
    po6676, po6677, po6678, po6679, po6680, po6681, po6682, po6683, po6684,
    po6685, po6686, po6687, po6688, po6689, po6690, po6691, po6692, po6693,
    po6694, po6695, po6696, po6697, po6698, po6699, po6700, po6701, po6702,
    po6703, po6704, po6705, po6706, po6707, po6708, po6709, po6710, po6711,
    po6712, po6713, po6714, po6715, po6716, po6717, po6718, po6719, po6720,
    po6721, po6722, po6723, po6724, po6725, po6726, po6727, po6728, po6729,
    po6730, po6731, po6732, po6733, po6734, po6735, po6736, po6737, po6738,
    po6739, po6740, po6741, po6742, po6743, po6744, po6745, po6746, po6747,
    po6748, po6749, po6750, po6751, po6752, po6753, po6754, po6755, po6756,
    po6757, po6758, po6759, po6760, po6761, po6762, po6763, po6764, po6765,
    po6766, po6767, po6768, po6769, po6770, po6771, po6772, po6773, po6774,
    po6775, po6776, po6777, po6778, po6779, po6780, po6781, po6782, po6783,
    po6784, po6785, po6786, po6787, po6788, po6789, po6790, po6791, po6792,
    po6793, po6794, po6795, po6796, po6797, po6798, po6799, po6800, po6801,
    po6802, po6803, po6804, po6805, po6806, po6807, po6808, po6809, po6810,
    po6811, po6812, po6813, po6814, po6815, po6816, po6817, po6818, po6819,
    po6820, po6821, po6822, po6823, po6824, po6825, po6826, po6827, po6828,
    po6829, po6830, po6831, po6832, po6833, po6834, po6835, po6836, po6837,
    po6838, po6839, po6840, po6841, po6842, po6843, po6844, po6845, po6846,
    po6847, po6848, po6849, po6850, po6851, po6852, po6853, po6854, po6855,
    po6856, po6857, po6858, po6859, po6860, po6861, po6862, po6863, po6864,
    po6865, po6866, po6867, po6868, po6869, po6870, po6871, po6872, po6873,
    po6874, po6875, po6876, po6877, po6878, po6879, po6880, po6881, po6882,
    po6883, po6884, po6885, po6886, po6887, po6888, po6889, po6890, po6891,
    po6892, po6893, po6894, po6895, po6896, po6897, po6898, po6899, po6900,
    po6901, po6902, po6903, po6904, po6905, po6906, po6907, po6908, po6909,
    po6910, po6911, po6912, po6913, po6914, po6915, po6916, po6917, po6918,
    po6919, po6920, po6921, po6922, po6923, po6924, po6925, po6926, po6927,
    po6928, po6929, po6930, po6931, po6932, po6933, po6934, po6935, po6936,
    po6937, po6938, po6939, po6940, po6941, po6942, po6943, po6944, po6945,
    po6946, po6947, po6948, po6949, po6950, po6951, po6952, po6953, po6954,
    po6955, po6956, po6957, po6958, po6959, po6960, po6961, po6962, po6963,
    po6964, po6965, po6966, po6967, po6968, po6969, po6970, po6971, po6972,
    po6973, po6974, po6975, po6976, po6977, po6978, po6979, po6980, po6981,
    po6982, po6983, po6984, po6985, po6986, po6987, po6988, po6989, po6990,
    po6991, po6992, po6993, po6994, po6995, po6996, po6997, po6998, po6999,
    po7000, po7001, po7002, po7003, po7004, po7005, po7006, po7007, po7008,
    po7009, po7010, po7011, po7012, po7013, po7014, po7015, po7016, po7017,
    po7018, po7019, po7020, po7021, po7022, po7023, po7024, po7025, po7026,
    po7027, po7028, po7029, po7030, po7031, po7032, po7033, po7034, po7035,
    po7036, po7037, po7038, po7039, po7040, po7041, po7042, po7043, po7044,
    po7045, po7046, po7047, po7048, po7049, po7050, po7051, po7052, po7053,
    po7054, po7055, po7056, po7057, po7058, po7059, po7060, po7061, po7062,
    po7063, po7064, po7065, po7066, po7067, po7068, po7069, po7070, po7071,
    po7072, po7073, po7074, po7075, po7076, po7077, po7078, po7079, po7080,
    po7081, po7082, po7083, po7084, po7085, po7086, po7087, po7088, po7089,
    po7090, po7091, po7092, po7093, po7094, po7095, po7096, po7097, po7098,
    po7099, po7100, po7101, po7102, po7103, po7104, po7105, po7106, po7107,
    po7108, po7109, po7110, po7111, po7112, po7113, po7114, po7115, po7116,
    po7117, po7118, po7119, po7120, po7121, po7122, po7123, po7124, po7125,
    po7126, po7127, po7128, po7129, po7130, po7131, po7132, po7133, po7134,
    po7135, po7136, po7137, po7138, po7139, po7140, po7141, po7142, po7143,
    po7144, po7145, po7146, po7147, po7148, po7149, po7150, po7151, po7152,
    po7153, po7154, po7155, po7156, po7157, po7158, po7159, po7160, po7161,
    po7162, po7163, po7164, po7165  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
    n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72,
    po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84,
    po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96,
    po97, po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125, po126,
    po127, po128, po129, po130, po131, po132, po133, po134, po135, po136,
    po137, po138, po139, po140, po141, po142, po143, po144, po145, po146,
    po147, po148, po149, po150, po151, po152, po153, po154, po155, po156,
    po157, po158, po159, po160, po161, po162, po163, po164, po165, po166,
    po167, po168, po169, po170, po171, po172, po173, po174, po175, po176,
    po177, po178, po179, po180, po181, po182, po183, po184, po185, po186,
    po187, po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215, po216,
    po217, po218, po219, po220, po221, po222, po223, po224, po225, po226,
    po227, po228, po229, po230, po231, po232, po233, po234, po235, po236,
    po237, po238, po239, po240, po241, po242, po243, po244, po245, po246,
    po247, po248, po249, po250, po251, po252, po253, po254, po255, po256,
    po257, po258, po259, po260, po261, po262, po263, po264, po265, po266,
    po267, po268, po269, po270, po271, po272, po273, po274, po275, po276,
    po277, po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305, po306,
    po307, po308, po309, po310, po311, po312, po313, po314, po315, po316,
    po317, po318, po319, po320, po321, po322, po323, po324, po325, po326,
    po327, po328, po329, po330, po331, po332, po333, po334, po335, po336,
    po337, po338, po339, po340, po341, po342, po343, po344, po345, po346,
    po347, po348, po349, po350, po351, po352, po353, po354, po355, po356,
    po357, po358, po359, po360, po361, po362, po363, po364, po365, po366,
    po367, po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395, po396,
    po397, po398, po399, po400, po401, po402, po403, po404, po405, po406,
    po407, po408, po409, po410, po411, po412, po413, po414, po415, po416,
    po417, po418, po419, po420, po421, po422, po423, po424, po425, po426,
    po427, po428, po429, po430, po431, po432, po433, po434, po435, po436,
    po437, po438, po439, po440, po441, po442, po443, po444, po445, po446,
    po447, po448, po449, po450, po451, po452, po453, po454, po455, po456,
    po457, po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485, po486,
    po487, po488, po489, po490, po491, po492, po493, po494, po495, po496,
    po497, po498, po499, po500, po501, po502, po503, po504, po505, po506,
    po507, po508, po509, po510, po511, po512, po513, po514, po515, po516,
    po517, po518, po519, po520, po521, po522, po523, po524, po525, po526,
    po527, po528, po529, po530, po531, po532, po533, po534, po535, po536,
    po537, po538, po539, po540, po541, po542, po543, po544, po545, po546,
    po547, po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575, po576,
    po577, po578, po579, po580, po581, po582, po583, po584, po585, po586,
    po587, po588, po589, po590, po591, po592, po593, po594, po595, po596,
    po597, po598, po599, po600, po601, po602, po603, po604, po605, po606,
    po607, po608, po609, po610, po611, po612, po613, po614, po615, po616,
    po617, po618, po619, po620, po621, po622, po623, po624, po625, po626,
    po627, po628, po629, po630, po631, po632, po633, po634, po635, po636,
    po637, po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665, po666,
    po667, po668, po669, po670, po671, po672, po673, po674, po675, po676,
    po677, po678, po679, po680, po681, po682, po683, po684, po685, po686,
    po687, po688, po689, po690, po691, po692, po693, po694, po695, po696,
    po697, po698, po699, po700, po701, po702, po703, po704, po705, po706,
    po707, po708, po709, po710, po711, po712, po713, po714, po715, po716,
    po717, po718, po719, po720, po721, po722, po723, po724, po725, po726,
    po727, po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755, po756,
    po757, po758, po759, po760, po761, po762, po763, po764, po765, po766,
    po767, po768, po769, po770, po771, po772, po773, po774, po775, po776,
    po777, po778, po779, po780, po781, po782, po783, po784, po785, po786,
    po787, po788, po789, po790, po791, po792, po793, po794, po795, po796,
    po797, po798, po799, po800, po801, po802, po803, po804, po805, po806,
    po807, po808, po809, po810, po811, po812, po813, po814, po815, po816,
    po817, po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845, po846,
    po847, po848, po849, po850, po851, po852, po853, po854, po855, po856,
    po857, po858, po859, po860, po861, po862, po863, po864, po865, po866,
    po867, po868, po869, po870, po871, po872, po873, po874, po875, po876,
    po877, po878, po879, po880, po881, po882, po883, po884, po885, po886,
    po887, po888, po889, po890, po891, po892, po893, po894, po895, po896,
    po897, po898, po899, po900, po901, po902, po903, po904, po905, po906,
    po907, po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935, po936,
    po937, po938, po939, po940, po941, po942, po943, po944, po945, po946,
    po947, po948, po949, po950, po951, po952, po953, po954, po955, po956,
    po957, po958, po959, po960, po961, po962, po963, po964, po965, po966,
    po967, po968, po969, po970, po971, po972, po973, po974, po975, po976,
    po977, po978, po979, po980, po981, po982, po983, po984, po985, po986,
    po987, po988, po989, po990, po991, po992, po993, po994, po995, po996,
    po997, po998, po999, po1000, po1001, po1002, po1003, po1004, po1005,
    po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014,
    po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023,
    po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032,
    po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041,
    po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050,
    po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059,
    po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068,
    po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077,
    po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086,
    po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095,
    po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104,
    po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113,
    po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122,
    po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131,
    po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140,
    po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149,
    po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158,
    po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167,
    po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176,
    po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185,
    po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194,
    po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203,
    po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212,
    po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221,
    po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230,
    po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239,
    po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248,
    po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257,
    po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266,
    po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275,
    po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284,
    po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293,
    po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302,
    po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311,
    po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320,
    po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329,
    po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338,
    po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347,
    po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356,
    po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365,
    po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374,
    po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383,
    po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392,
    po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401,
    po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410,
    po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419,
    po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428,
    po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437,
    po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446,
    po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455,
    po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464,
    po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473,
    po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482,
    po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491,
    po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500,
    po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509,
    po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518,
    po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527,
    po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536,
    po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545,
    po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554,
    po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563,
    po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572,
    po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581,
    po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590,
    po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599,
    po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608,
    po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617,
    po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626,
    po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635,
    po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644,
    po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653,
    po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662,
    po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671,
    po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680,
    po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689,
    po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698,
    po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707,
    po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716,
    po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725,
    po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734,
    po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743,
    po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752,
    po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761,
    po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770,
    po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779,
    po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788,
    po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797,
    po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806,
    po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815,
    po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824,
    po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833,
    po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842,
    po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851,
    po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860,
    po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869,
    po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878,
    po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887,
    po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896,
    po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905,
    po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914,
    po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923,
    po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932,
    po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941,
    po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950,
    po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959,
    po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968,
    po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977,
    po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986,
    po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995,
    po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004,
    po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013,
    po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022,
    po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031,
    po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040,
    po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049,
    po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058,
    po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067,
    po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076,
    po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085,
    po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094,
    po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103,
    po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112,
    po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121,
    po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130,
    po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139,
    po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148,
    po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157,
    po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166,
    po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175,
    po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184,
    po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193,
    po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202,
    po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211,
    po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220,
    po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229,
    po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238,
    po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247,
    po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256,
    po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265,
    po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274,
    po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283,
    po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292,
    po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301,
    po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310,
    po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319,
    po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328,
    po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337,
    po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346,
    po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355,
    po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364,
    po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373,
    po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382,
    po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391,
    po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400,
    po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409,
    po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418,
    po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427,
    po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436,
    po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445,
    po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454,
    po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463,
    po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472,
    po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481,
    po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490,
    po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499,
    po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508,
    po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517,
    po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526,
    po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535,
    po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544,
    po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553,
    po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562,
    po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571,
    po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580,
    po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589,
    po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598,
    po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607,
    po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616,
    po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625,
    po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634,
    po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643,
    po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652,
    po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661,
    po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670,
    po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679,
    po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688,
    po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697,
    po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706,
    po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715,
    po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724,
    po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733,
    po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742,
    po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751,
    po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760,
    po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769,
    po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778,
    po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787,
    po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796,
    po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805,
    po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814,
    po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823,
    po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832,
    po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841,
    po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850,
    po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859,
    po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868,
    po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877,
    po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886,
    po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895,
    po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904,
    po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913,
    po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922,
    po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931,
    po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940,
    po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949,
    po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958,
    po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967,
    po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976,
    po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985,
    po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994,
    po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003,
    po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012,
    po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021,
    po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030,
    po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039,
    po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048,
    po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057,
    po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066,
    po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075,
    po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084,
    po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093,
    po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102,
    po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111,
    po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120,
    po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129,
    po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138,
    po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147,
    po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156,
    po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165,
    po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174,
    po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183,
    po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192,
    po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201,
    po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210,
    po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219,
    po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228,
    po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237,
    po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246,
    po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255,
    po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264,
    po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273,
    po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282,
    po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291,
    po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300,
    po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309,
    po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318,
    po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327,
    po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336,
    po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345,
    po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354,
    po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363,
    po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372,
    po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381,
    po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390,
    po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399,
    po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408,
    po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417,
    po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426,
    po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435,
    po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444,
    po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453,
    po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462,
    po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471,
    po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480,
    po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489,
    po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498,
    po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507,
    po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516,
    po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525,
    po3526, po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534,
    po3535, po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543,
    po3544, po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552,
    po3553, po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561,
    po3562, po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570,
    po3571, po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579,
    po3580, po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588,
    po3589, po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597,
    po3598, po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606,
    po3607, po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615,
    po3616, po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624,
    po3625, po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633,
    po3634, po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642,
    po3643, po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651,
    po3652, po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660,
    po3661, po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669,
    po3670, po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678,
    po3679, po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687,
    po3688, po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696,
    po3697, po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705,
    po3706, po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714,
    po3715, po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723,
    po3724, po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732,
    po3733, po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741,
    po3742, po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750,
    po3751, po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759,
    po3760, po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768,
    po3769, po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777,
    po3778, po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786,
    po3787, po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795,
    po3796, po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804,
    po3805, po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813,
    po3814, po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822,
    po3823, po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831,
    po3832, po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840,
    po3841, po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849,
    po3850, po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858,
    po3859, po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867,
    po3868, po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876,
    po3877, po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885,
    po3886, po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894,
    po3895, po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903,
    po3904, po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912,
    po3913, po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921,
    po3922, po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930,
    po3931, po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939,
    po3940, po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948,
    po3949, po3950, po3951, po3952, po3953, po3954, po3955, po3956, po3957,
    po3958, po3959, po3960, po3961, po3962, po3963, po3964, po3965, po3966,
    po3967, po3968, po3969, po3970, po3971, po3972, po3973, po3974, po3975,
    po3976, po3977, po3978, po3979, po3980, po3981, po3982, po3983, po3984,
    po3985, po3986, po3987, po3988, po3989, po3990, po3991, po3992, po3993,
    po3994, po3995, po3996, po3997, po3998, po3999, po4000, po4001, po4002,
    po4003, po4004, po4005, po4006, po4007, po4008, po4009, po4010, po4011,
    po4012, po4013, po4014, po4015, po4016, po4017, po4018, po4019, po4020,
    po4021, po4022, po4023, po4024, po4025, po4026, po4027, po4028, po4029,
    po4030, po4031, po4032, po4033, po4034, po4035, po4036, po4037, po4038,
    po4039, po4040, po4041, po4042, po4043, po4044, po4045, po4046, po4047,
    po4048, po4049, po4050, po4051, po4052, po4053, po4054, po4055, po4056,
    po4057, po4058, po4059, po4060, po4061, po4062, po4063, po4064, po4065,
    po4066, po4067, po4068, po4069, po4070, po4071, po4072, po4073, po4074,
    po4075, po4076, po4077, po4078, po4079, po4080, po4081, po4082, po4083,
    po4084, po4085, po4086, po4087, po4088, po4089, po4090, po4091, po4092,
    po4093, po4094, po4095, po4096, po4097, po4098, po4099, po4100, po4101,
    po4102, po4103, po4104, po4105, po4106, po4107, po4108, po4109, po4110,
    po4111, po4112, po4113, po4114, po4115, po4116, po4117, po4118, po4119,
    po4120, po4121, po4122, po4123, po4124, po4125, po4126, po4127, po4128,
    po4129, po4130, po4131, po4132, po4133, po4134, po4135, po4136, po4137,
    po4138, po4139, po4140, po4141, po4142, po4143, po4144, po4145, po4146,
    po4147, po4148, po4149, po4150, po4151, po4152, po4153, po4154, po4155,
    po4156, po4157, po4158, po4159, po4160, po4161, po4162, po4163, po4164,
    po4165, po4166, po4167, po4168, po4169, po4170, po4171, po4172, po4173,
    po4174, po4175, po4176, po4177, po4178, po4179, po4180, po4181, po4182,
    po4183, po4184, po4185, po4186, po4187, po4188, po4189, po4190, po4191,
    po4192, po4193, po4194, po4195, po4196, po4197, po4198, po4199, po4200,
    po4201, po4202, po4203, po4204, po4205, po4206, po4207, po4208, po4209,
    po4210, po4211, po4212, po4213, po4214, po4215, po4216, po4217, po4218,
    po4219, po4220, po4221, po4222, po4223, po4224, po4225, po4226, po4227,
    po4228, po4229, po4230, po4231, po4232, po4233, po4234, po4235, po4236,
    po4237, po4238, po4239, po4240, po4241, po4242, po4243, po4244, po4245,
    po4246, po4247, po4248, po4249, po4250, po4251, po4252, po4253, po4254,
    po4255, po4256, po4257, po4258, po4259, po4260, po4261, po4262, po4263,
    po4264, po4265, po4266, po4267, po4268, po4269, po4270, po4271, po4272,
    po4273, po4274, po4275, po4276, po4277, po4278, po4279, po4280, po4281,
    po4282, po4283, po4284, po4285, po4286, po4287, po4288, po4289, po4290,
    po4291, po4292, po4293, po4294, po4295, po4296, po4297, po4298, po4299,
    po4300, po4301, po4302, po4303, po4304, po4305, po4306, po4307, po4308,
    po4309, po4310, po4311, po4312, po4313, po4314, po4315, po4316, po4317,
    po4318, po4319, po4320, po4321, po4322, po4323, po4324, po4325, po4326,
    po4327, po4328, po4329, po4330, po4331, po4332, po4333, po4334, po4335,
    po4336, po4337, po4338, po4339, po4340, po4341, po4342, po4343, po4344,
    po4345, po4346, po4347, po4348, po4349, po4350, po4351, po4352, po4353,
    po4354, po4355, po4356, po4357, po4358, po4359, po4360, po4361, po4362,
    po4363, po4364, po4365, po4366, po4367, po4368, po4369, po4370, po4371,
    po4372, po4373, po4374, po4375, po4376, po4377, po4378, po4379, po4380,
    po4381, po4382, po4383, po4384, po4385, po4386, po4387, po4388, po4389,
    po4390, po4391, po4392, po4393, po4394, po4395, po4396, po4397, po4398,
    po4399, po4400, po4401, po4402, po4403, po4404, po4405, po4406, po4407,
    po4408, po4409, po4410, po4411, po4412, po4413, po4414, po4415, po4416,
    po4417, po4418, po4419, po4420, po4421, po4422, po4423, po4424, po4425,
    po4426, po4427, po4428, po4429, po4430, po4431, po4432, po4433, po4434,
    po4435, po4436, po4437, po4438, po4439, po4440, po4441, po4442, po4443,
    po4444, po4445, po4446, po4447, po4448, po4449, po4450, po4451, po4452,
    po4453, po4454, po4455, po4456, po4457, po4458, po4459, po4460, po4461,
    po4462, po4463, po4464, po4465, po4466, po4467, po4468, po4469, po4470,
    po4471, po4472, po4473, po4474, po4475, po4476, po4477, po4478, po4479,
    po4480, po4481, po4482, po4483, po4484, po4485, po4486, po4487, po4488,
    po4489, po4490, po4491, po4492, po4493, po4494, po4495, po4496, po4497,
    po4498, po4499, po4500, po4501, po4502, po4503, po4504, po4505, po4506,
    po4507, po4508, po4509, po4510, po4511, po4512, po4513, po4514, po4515,
    po4516, po4517, po4518, po4519, po4520, po4521, po4522, po4523, po4524,
    po4525, po4526, po4527, po4528, po4529, po4530, po4531, po4532, po4533,
    po4534, po4535, po4536, po4537, po4538, po4539, po4540, po4541, po4542,
    po4543, po4544, po4545, po4546, po4547, po4548, po4549, po4550, po4551,
    po4552, po4553, po4554, po4555, po4556, po4557, po4558, po4559, po4560,
    po4561, po4562, po4563, po4564, po4565, po4566, po4567, po4568, po4569,
    po4570, po4571, po4572, po4573, po4574, po4575, po4576, po4577, po4578,
    po4579, po4580, po4581, po4582, po4583, po4584, po4585, po4586, po4587,
    po4588, po4589, po4590, po4591, po4592, po4593, po4594, po4595, po4596,
    po4597, po4598, po4599, po4600, po4601, po4602, po4603, po4604, po4605,
    po4606, po4607, po4608, po4609, po4610, po4611, po4612, po4613, po4614,
    po4615, po4616, po4617, po4618, po4619, po4620, po4621, po4622, po4623,
    po4624, po4625, po4626, po4627, po4628, po4629, po4630, po4631, po4632,
    po4633, po4634, po4635, po4636, po4637, po4638, po4639, po4640, po4641,
    po4642, po4643, po4644, po4645, po4646, po4647, po4648, po4649, po4650,
    po4651, po4652, po4653, po4654, po4655, po4656, po4657, po4658, po4659,
    po4660, po4661, po4662, po4663, po4664, po4665, po4666, po4667, po4668,
    po4669, po4670, po4671, po4672, po4673, po4674, po4675, po4676, po4677,
    po4678, po4679, po4680, po4681, po4682, po4683, po4684, po4685, po4686,
    po4687, po4688, po4689, po4690, po4691, po4692, po4693, po4694, po4695,
    po4696, po4697, po4698, po4699, po4700, po4701, po4702, po4703, po4704,
    po4705, po4706, po4707, po4708, po4709, po4710, po4711, po4712, po4713,
    po4714, po4715, po4716, po4717, po4718, po4719, po4720, po4721, po4722,
    po4723, po4724, po4725, po4726, po4727, po4728, po4729, po4730, po4731,
    po4732, po4733, po4734, po4735, po4736, po4737, po4738, po4739, po4740,
    po4741, po4742, po4743, po4744, po4745, po4746, po4747, po4748, po4749,
    po4750, po4751, po4752, po4753, po4754, po4755, po4756, po4757, po4758,
    po4759, po4760, po4761, po4762, po4763, po4764, po4765, po4766, po4767,
    po4768, po4769, po4770, po4771, po4772, po4773, po4774, po4775, po4776,
    po4777, po4778, po4779, po4780, po4781, po4782, po4783, po4784, po4785,
    po4786, po4787, po4788, po4789, po4790, po4791, po4792, po4793, po4794,
    po4795, po4796, po4797, po4798, po4799, po4800, po4801, po4802, po4803,
    po4804, po4805, po4806, po4807, po4808, po4809, po4810, po4811, po4812,
    po4813, po4814, po4815, po4816, po4817, po4818, po4819, po4820, po4821,
    po4822, po4823, po4824, po4825, po4826, po4827, po4828, po4829, po4830,
    po4831, po4832, po4833, po4834, po4835, po4836, po4837, po4838, po4839,
    po4840, po4841, po4842, po4843, po4844, po4845, po4846, po4847, po4848,
    po4849, po4850, po4851, po4852, po4853, po4854, po4855, po4856, po4857,
    po4858, po4859, po4860, po4861, po4862, po4863, po4864, po4865, po4866,
    po4867, po4868, po4869, po4870, po4871, po4872, po4873, po4874, po4875,
    po4876, po4877, po4878, po4879, po4880, po4881, po4882, po4883, po4884,
    po4885, po4886, po4887, po4888, po4889, po4890, po4891, po4892, po4893,
    po4894, po4895, po4896, po4897, po4898, po4899, po4900, po4901, po4902,
    po4903, po4904, po4905, po4906, po4907, po4908, po4909, po4910, po4911,
    po4912, po4913, po4914, po4915, po4916, po4917, po4918, po4919, po4920,
    po4921, po4922, po4923, po4924, po4925, po4926, po4927, po4928, po4929,
    po4930, po4931, po4932, po4933, po4934, po4935, po4936, po4937, po4938,
    po4939, po4940, po4941, po4942, po4943, po4944, po4945, po4946, po4947,
    po4948, po4949, po4950, po4951, po4952, po4953, po4954, po4955, po4956,
    po4957, po4958, po4959, po4960, po4961, po4962, po4963, po4964, po4965,
    po4966, po4967, po4968, po4969, po4970, po4971, po4972, po4973, po4974,
    po4975, po4976, po4977, po4978, po4979, po4980, po4981, po4982, po4983,
    po4984, po4985, po4986, po4987, po4988, po4989, po4990, po4991, po4992,
    po4993, po4994, po4995, po4996, po4997, po4998, po4999, po5000, po5001,
    po5002, po5003, po5004, po5005, po5006, po5007, po5008, po5009, po5010,
    po5011, po5012, po5013, po5014, po5015, po5016, po5017, po5018, po5019,
    po5020, po5021, po5022, po5023, po5024, po5025, po5026, po5027, po5028,
    po5029, po5030, po5031, po5032, po5033, po5034, po5035, po5036, po5037,
    po5038, po5039, po5040, po5041, po5042, po5043, po5044, po5045, po5046,
    po5047, po5048, po5049, po5050, po5051, po5052, po5053, po5054, po5055,
    po5056, po5057, po5058, po5059, po5060, po5061, po5062, po5063, po5064,
    po5065, po5066, po5067, po5068, po5069, po5070, po5071, po5072, po5073,
    po5074, po5075, po5076, po5077, po5078, po5079, po5080, po5081, po5082,
    po5083, po5084, po5085, po5086, po5087, po5088, po5089, po5090, po5091,
    po5092, po5093, po5094, po5095, po5096, po5097, po5098, po5099, po5100,
    po5101, po5102, po5103, po5104, po5105, po5106, po5107, po5108, po5109,
    po5110, po5111, po5112, po5113, po5114, po5115, po5116, po5117, po5118,
    po5119, po5120, po5121, po5122, po5123, po5124, po5125, po5126, po5127,
    po5128, po5129, po5130, po5131, po5132, po5133, po5134, po5135, po5136,
    po5137, po5138, po5139, po5140, po5141, po5142, po5143, po5144, po5145,
    po5146, po5147, po5148, po5149, po5150, po5151, po5152, po5153, po5154,
    po5155, po5156, po5157, po5158, po5159, po5160, po5161, po5162, po5163,
    po5164, po5165, po5166, po5167, po5168, po5169, po5170, po5171, po5172,
    po5173, po5174, po5175, po5176, po5177, po5178, po5179, po5180, po5181,
    po5182, po5183, po5184, po5185, po5186, po5187, po5188, po5189, po5190,
    po5191, po5192, po5193, po5194, po5195, po5196, po5197, po5198, po5199,
    po5200, po5201, po5202, po5203, po5204, po5205, po5206, po5207, po5208,
    po5209, po5210, po5211, po5212, po5213, po5214, po5215, po5216, po5217,
    po5218, po5219, po5220, po5221, po5222, po5223, po5224, po5225, po5226,
    po5227, po5228, po5229, po5230, po5231, po5232, po5233, po5234, po5235,
    po5236, po5237, po5238, po5239, po5240, po5241, po5242, po5243, po5244,
    po5245, po5246, po5247, po5248, po5249, po5250, po5251, po5252, po5253,
    po5254, po5255, po5256, po5257, po5258, po5259, po5260, po5261, po5262,
    po5263, po5264, po5265, po5266, po5267, po5268, po5269, po5270, po5271,
    po5272, po5273, po5274, po5275, po5276, po5277, po5278, po5279, po5280,
    po5281, po5282, po5283, po5284, po5285, po5286, po5287, po5288, po5289,
    po5290, po5291, po5292, po5293, po5294, po5295, po5296, po5297, po5298,
    po5299, po5300, po5301, po5302, po5303, po5304, po5305, po5306, po5307,
    po5308, po5309, po5310, po5311, po5312, po5313, po5314, po5315, po5316,
    po5317, po5318, po5319, po5320, po5321, po5322, po5323, po5324, po5325,
    po5326, po5327, po5328, po5329, po5330, po5331, po5332, po5333, po5334,
    po5335, po5336, po5337, po5338, po5339, po5340, po5341, po5342, po5343,
    po5344, po5345, po5346, po5347, po5348, po5349, po5350, po5351, po5352,
    po5353, po5354, po5355, po5356, po5357, po5358, po5359, po5360, po5361,
    po5362, po5363, po5364, po5365, po5366, po5367, po5368, po5369, po5370,
    po5371, po5372, po5373, po5374, po5375, po5376, po5377, po5378, po5379,
    po5380, po5381, po5382, po5383, po5384, po5385, po5386, po5387, po5388,
    po5389, po5390, po5391, po5392, po5393, po5394, po5395, po5396, po5397,
    po5398, po5399, po5400, po5401, po5402, po5403, po5404, po5405, po5406,
    po5407, po5408, po5409, po5410, po5411, po5412, po5413, po5414, po5415,
    po5416, po5417, po5418, po5419, po5420, po5421, po5422, po5423, po5424,
    po5425, po5426, po5427, po5428, po5429, po5430, po5431, po5432, po5433,
    po5434, po5435, po5436, po5437, po5438, po5439, po5440, po5441, po5442,
    po5443, po5444, po5445, po5446, po5447, po5448, po5449, po5450, po5451,
    po5452, po5453, po5454, po5455, po5456, po5457, po5458, po5459, po5460,
    po5461, po5462, po5463, po5464, po5465, po5466, po5467, po5468, po5469,
    po5470, po5471, po5472, po5473, po5474, po5475, po5476, po5477, po5478,
    po5479, po5480, po5481, po5482, po5483, po5484, po5485, po5486, po5487,
    po5488, po5489, po5490, po5491, po5492, po5493, po5494, po5495, po5496,
    po5497, po5498, po5499, po5500, po5501, po5502, po5503, po5504, po5505,
    po5506, po5507, po5508, po5509, po5510, po5511, po5512, po5513, po5514,
    po5515, po5516, po5517, po5518, po5519, po5520, po5521, po5522, po5523,
    po5524, po5525, po5526, po5527, po5528, po5529, po5530, po5531, po5532,
    po5533, po5534, po5535, po5536, po5537, po5538, po5539, po5540, po5541,
    po5542, po5543, po5544, po5545, po5546, po5547, po5548, po5549, po5550,
    po5551, po5552, po5553, po5554, po5555, po5556, po5557, po5558, po5559,
    po5560, po5561, po5562, po5563, po5564, po5565, po5566, po5567, po5568,
    po5569, po5570, po5571, po5572, po5573, po5574, po5575, po5576, po5577,
    po5578, po5579, po5580, po5581, po5582, po5583, po5584, po5585, po5586,
    po5587, po5588, po5589, po5590, po5591, po5592, po5593, po5594, po5595,
    po5596, po5597, po5598, po5599, po5600, po5601, po5602, po5603, po5604,
    po5605, po5606, po5607, po5608, po5609, po5610, po5611, po5612, po5613,
    po5614, po5615, po5616, po5617, po5618, po5619, po5620, po5621, po5622,
    po5623, po5624, po5625, po5626, po5627, po5628, po5629, po5630, po5631,
    po5632, po5633, po5634, po5635, po5636, po5637, po5638, po5639, po5640,
    po5641, po5642, po5643, po5644, po5645, po5646, po5647, po5648, po5649,
    po5650, po5651, po5652, po5653, po5654, po5655, po5656, po5657, po5658,
    po5659, po5660, po5661, po5662, po5663, po5664, po5665, po5666, po5667,
    po5668, po5669, po5670, po5671, po5672, po5673, po5674, po5675, po5676,
    po5677, po5678, po5679, po5680, po5681, po5682, po5683, po5684, po5685,
    po5686, po5687, po5688, po5689, po5690, po5691, po5692, po5693, po5694,
    po5695, po5696, po5697, po5698, po5699, po5700, po5701, po5702, po5703,
    po5704, po5705, po5706, po5707, po5708, po5709, po5710, po5711, po5712,
    po5713, po5714, po5715, po5716, po5717, po5718, po5719, po5720, po5721,
    po5722, po5723, po5724, po5725, po5726, po5727, po5728, po5729, po5730,
    po5731, po5732, po5733, po5734, po5735, po5736, po5737, po5738, po5739,
    po5740, po5741, po5742, po5743, po5744, po5745, po5746, po5747, po5748,
    po5749, po5750, po5751, po5752, po5753, po5754, po5755, po5756, po5757,
    po5758, po5759, po5760, po5761, po5762, po5763, po5764, po5765, po5766,
    po5767, po5768, po5769, po5770, po5771, po5772, po5773, po5774, po5775,
    po5776, po5777, po5778, po5779, po5780, po5781, po5782, po5783, po5784,
    po5785, po5786, po5787, po5788, po5789, po5790, po5791, po5792, po5793,
    po5794, po5795, po5796, po5797, po5798, po5799, po5800, po5801, po5802,
    po5803, po5804, po5805, po5806, po5807, po5808, po5809, po5810, po5811,
    po5812, po5813, po5814, po5815, po5816, po5817, po5818, po5819, po5820,
    po5821, po5822, po5823, po5824, po5825, po5826, po5827, po5828, po5829,
    po5830, po5831, po5832, po5833, po5834, po5835, po5836, po5837, po5838,
    po5839, po5840, po5841, po5842, po5843, po5844, po5845, po5846, po5847,
    po5848, po5849, po5850, po5851, po5852, po5853, po5854, po5855, po5856,
    po5857, po5858, po5859, po5860, po5861, po5862, po5863, po5864, po5865,
    po5866, po5867, po5868, po5869, po5870, po5871, po5872, po5873, po5874,
    po5875, po5876, po5877, po5878, po5879, po5880, po5881, po5882, po5883,
    po5884, po5885, po5886, po5887, po5888, po5889, po5890, po5891, po5892,
    po5893, po5894, po5895, po5896, po5897, po5898, po5899, po5900, po5901,
    po5902, po5903, po5904, po5905, po5906, po5907, po5908, po5909, po5910,
    po5911, po5912, po5913, po5914, po5915, po5916, po5917, po5918, po5919,
    po5920, po5921, po5922, po5923, po5924, po5925, po5926, po5927, po5928,
    po5929, po5930, po5931, po5932, po5933, po5934, po5935, po5936, po5937,
    po5938, po5939, po5940, po5941, po5942, po5943, po5944, po5945, po5946,
    po5947, po5948, po5949, po5950, po5951, po5952, po5953, po5954, po5955,
    po5956, po5957, po5958, po5959, po5960, po5961, po5962, po5963, po5964,
    po5965, po5966, po5967, po5968, po5969, po5970, po5971, po5972, po5973,
    po5974, po5975, po5976, po5977, po5978, po5979, po5980, po5981, po5982,
    po5983, po5984, po5985, po5986, po5987, po5988, po5989, po5990, po5991,
    po5992, po5993, po5994, po5995, po5996, po5997, po5998, po5999, po6000,
    po6001, po6002, po6003, po6004, po6005, po6006, po6007, po6008, po6009,
    po6010, po6011, po6012, po6013, po6014, po6015, po6016, po6017, po6018,
    po6019, po6020, po6021, po6022, po6023, po6024, po6025, po6026, po6027,
    po6028, po6029, po6030, po6031, po6032, po6033, po6034, po6035, po6036,
    po6037, po6038, po6039, po6040, po6041, po6042, po6043, po6044, po6045,
    po6046, po6047, po6048, po6049, po6050, po6051, po6052, po6053, po6054,
    po6055, po6056, po6057, po6058, po6059, po6060, po6061, po6062, po6063,
    po6064, po6065, po6066, po6067, po6068, po6069, po6070, po6071, po6072,
    po6073, po6074, po6075, po6076, po6077, po6078, po6079, po6080, po6081,
    po6082, po6083, po6084, po6085, po6086, po6087, po6088, po6089, po6090,
    po6091, po6092, po6093, po6094, po6095, po6096, po6097, po6098, po6099,
    po6100, po6101, po6102, po6103, po6104, po6105, po6106, po6107, po6108,
    po6109, po6110, po6111, po6112, po6113, po6114, po6115, po6116, po6117,
    po6118, po6119, po6120, po6121, po6122, po6123, po6124, po6125, po6126,
    po6127, po6128, po6129, po6130, po6131, po6132, po6133, po6134, po6135,
    po6136, po6137, po6138, po6139, po6140, po6141, po6142, po6143, po6144,
    po6145, po6146, po6147, po6148, po6149, po6150, po6151, po6152, po6153,
    po6154, po6155, po6156, po6157, po6158, po6159, po6160, po6161, po6162,
    po6163, po6164, po6165, po6166, po6167, po6168, po6169, po6170, po6171,
    po6172, po6173, po6174, po6175, po6176, po6177, po6178, po6179, po6180,
    po6181, po6182, po6183, po6184, po6185, po6186, po6187, po6188, po6189,
    po6190, po6191, po6192, po6193, po6194, po6195, po6196, po6197, po6198,
    po6199, po6200, po6201, po6202, po6203, po6204, po6205, po6206, po6207,
    po6208, po6209, po6210, po6211, po6212, po6213, po6214, po6215, po6216,
    po6217, po6218, po6219, po6220, po6221, po6222, po6223, po6224, po6225,
    po6226, po6227, po6228, po6229, po6230, po6231, po6232, po6233, po6234,
    po6235, po6236, po6237, po6238, po6239, po6240, po6241, po6242, po6243,
    po6244, po6245, po6246, po6247, po6248, po6249, po6250, po6251, po6252,
    po6253, po6254, po6255, po6256, po6257, po6258, po6259, po6260, po6261,
    po6262, po6263, po6264, po6265, po6266, po6267, po6268, po6269, po6270,
    po6271, po6272, po6273, po6274, po6275, po6276, po6277, po6278, po6279,
    po6280, po6281, po6282, po6283, po6284, po6285, po6286, po6287, po6288,
    po6289, po6290, po6291, po6292, po6293, po6294, po6295, po6296, po6297,
    po6298, po6299, po6300, po6301, po6302, po6303, po6304, po6305, po6306,
    po6307, po6308, po6309, po6310, po6311, po6312, po6313, po6314, po6315,
    po6316, po6317, po6318, po6319, po6320, po6321, po6322, po6323, po6324,
    po6325, po6326, po6327, po6328, po6329, po6330, po6331, po6332, po6333,
    po6334, po6335, po6336, po6337, po6338, po6339, po6340, po6341, po6342,
    po6343, po6344, po6345, po6346, po6347, po6348, po6349, po6350, po6351,
    po6352, po6353, po6354, po6355, po6356, po6357, po6358, po6359, po6360,
    po6361, po6362, po6363, po6364, po6365, po6366, po6367, po6368, po6369,
    po6370, po6371, po6372, po6373, po6374, po6375, po6376, po6377, po6378,
    po6379, po6380, po6381, po6382, po6383, po6384, po6385, po6386, po6387,
    po6388, po6389, po6390, po6391, po6392, po6393, po6394, po6395, po6396,
    po6397, po6398, po6399, po6400, po6401, po6402, po6403, po6404, po6405,
    po6406, po6407, po6408, po6409, po6410, po6411, po6412, po6413, po6414,
    po6415, po6416, po6417, po6418, po6419, po6420, po6421, po6422, po6423,
    po6424, po6425, po6426, po6427, po6428, po6429, po6430, po6431, po6432,
    po6433, po6434, po6435, po6436, po6437, po6438, po6439, po6440, po6441,
    po6442, po6443, po6444, po6445, po6446, po6447, po6448, po6449, po6450,
    po6451, po6452, po6453, po6454, po6455, po6456, po6457, po6458, po6459,
    po6460, po6461, po6462, po6463, po6464, po6465, po6466, po6467, po6468,
    po6469, po6470, po6471, po6472, po6473, po6474, po6475, po6476, po6477,
    po6478, po6479, po6480, po6481, po6482, po6483, po6484, po6485, po6486,
    po6487, po6488, po6489, po6490, po6491, po6492, po6493, po6494, po6495,
    po6496, po6497, po6498, po6499, po6500, po6501, po6502, po6503, po6504,
    po6505, po6506, po6507, po6508, po6509, po6510, po6511, po6512, po6513,
    po6514, po6515, po6516, po6517, po6518, po6519, po6520, po6521, po6522,
    po6523, po6524, po6525, po6526, po6527, po6528, po6529, po6530, po6531,
    po6532, po6533, po6534, po6535, po6536, po6537, po6538, po6539, po6540,
    po6541, po6542, po6543, po6544, po6545, po6546, po6547, po6548, po6549,
    po6550, po6551, po6552, po6553, po6554, po6555, po6556, po6557, po6558,
    po6559, po6560, po6561, po6562, po6563, po6564, po6565, po6566, po6567,
    po6568, po6569, po6570, po6571, po6572, po6573, po6574, po6575, po6576,
    po6577, po6578, po6579, po6580, po6581, po6582, po6583, po6584, po6585,
    po6586, po6587, po6588, po6589, po6590, po6591, po6592, po6593, po6594,
    po6595, po6596, po6597, po6598, po6599, po6600, po6601, po6602, po6603,
    po6604, po6605, po6606, po6607, po6608, po6609, po6610, po6611, po6612,
    po6613, po6614, po6615, po6616, po6617, po6618, po6619, po6620, po6621,
    po6622, po6623, po6624, po6625, po6626, po6627, po6628, po6629, po6630,
    po6631, po6632, po6633, po6634, po6635, po6636, po6637, po6638, po6639,
    po6640, po6641, po6642, po6643, po6644, po6645, po6646, po6647, po6648,
    po6649, po6650, po6651, po6652, po6653, po6654, po6655, po6656, po6657,
    po6658, po6659, po6660, po6661, po6662, po6663, po6664, po6665, po6666,
    po6667, po6668, po6669, po6670, po6671, po6672, po6673, po6674, po6675,
    po6676, po6677, po6678, po6679, po6680, po6681, po6682, po6683, po6684,
    po6685, po6686, po6687, po6688, po6689, po6690, po6691, po6692, po6693,
    po6694, po6695, po6696, po6697, po6698, po6699, po6700, po6701, po6702,
    po6703, po6704, po6705, po6706, po6707, po6708, po6709, po6710, po6711,
    po6712, po6713, po6714, po6715, po6716, po6717, po6718, po6719, po6720,
    po6721, po6722, po6723, po6724, po6725, po6726, po6727, po6728, po6729,
    po6730, po6731, po6732, po6733, po6734, po6735, po6736, po6737, po6738,
    po6739, po6740, po6741, po6742, po6743, po6744, po6745, po6746, po6747,
    po6748, po6749, po6750, po6751, po6752, po6753, po6754, po6755, po6756,
    po6757, po6758, po6759, po6760, po6761, po6762, po6763, po6764, po6765,
    po6766, po6767, po6768, po6769, po6770, po6771, po6772, po6773, po6774,
    po6775, po6776, po6777, po6778, po6779, po6780, po6781, po6782, po6783,
    po6784, po6785, po6786, po6787, po6788, po6789, po6790, po6791, po6792,
    po6793, po6794, po6795, po6796, po6797, po6798, po6799, po6800, po6801,
    po6802, po6803, po6804, po6805, po6806, po6807, po6808, po6809, po6810,
    po6811, po6812, po6813, po6814, po6815, po6816, po6817, po6818, po6819,
    po6820, po6821, po6822, po6823, po6824, po6825, po6826, po6827, po6828,
    po6829, po6830, po6831, po6832, po6833, po6834, po6835, po6836, po6837,
    po6838, po6839, po6840, po6841, po6842, po6843, po6844, po6845, po6846,
    po6847, po6848, po6849, po6850, po6851, po6852, po6853, po6854, po6855,
    po6856, po6857, po6858, po6859, po6860, po6861, po6862, po6863, po6864,
    po6865, po6866, po6867, po6868, po6869, po6870, po6871, po6872, po6873,
    po6874, po6875, po6876, po6877, po6878, po6879, po6880, po6881, po6882,
    po6883, po6884, po6885, po6886, po6887, po6888, po6889, po6890, po6891,
    po6892, po6893, po6894, po6895, po6896, po6897, po6898, po6899, po6900,
    po6901, po6902, po6903, po6904, po6905, po6906, po6907, po6908, po6909,
    po6910, po6911, po6912, po6913, po6914, po6915, po6916, po6917, po6918,
    po6919, po6920, po6921, po6922, po6923, po6924, po6925, po6926, po6927,
    po6928, po6929, po6930, po6931, po6932, po6933, po6934, po6935, po6936,
    po6937, po6938, po6939, po6940, po6941, po6942, po6943, po6944, po6945,
    po6946, po6947, po6948, po6949, po6950, po6951, po6952, po6953, po6954,
    po6955, po6956, po6957, po6958, po6959, po6960, po6961, po6962, po6963,
    po6964, po6965, po6966, po6967, po6968, po6969, po6970, po6971, po6972,
    po6973, po6974, po6975, po6976, po6977, po6978, po6979, po6980, po6981,
    po6982, po6983, po6984, po6985, po6986, po6987, po6988, po6989, po6990,
    po6991, po6992, po6993, po6994, po6995, po6996, po6997, po6998, po6999,
    po7000, po7001, po7002, po7003, po7004, po7005, po7006, po7007, po7008,
    po7009, po7010, po7011, po7012, po7013, po7014, po7015, po7016, po7017,
    po7018, po7019, po7020, po7021, po7022, po7023, po7024, po7025, po7026,
    po7027, po7028, po7029, po7030, po7031, po7032, po7033, po7034, po7035,
    po7036, po7037, po7038, po7039, po7040, po7041, po7042, po7043, po7044,
    po7045, po7046, po7047, po7048, po7049, po7050, po7051, po7052, po7053,
    po7054, po7055, po7056, po7057, po7058, po7059, po7060, po7061, po7062,
    po7063, po7064, po7065, po7066, po7067, po7068, po7069, po7070, po7071,
    po7072, po7073, po7074, po7075, po7076, po7077, po7078, po7079, po7080,
    po7081, po7082, po7083, po7084, po7085, po7086, po7087, po7088, po7089,
    po7090, po7091, po7092, po7093, po7094, po7095, po7096, po7097, po7098,
    po7099, po7100, po7101, po7102, po7103, po7104, po7105, po7106, po7107,
    po7108, po7109, po7110, po7111, po7112, po7113, po7114, po7115, po7116,
    po7117, po7118, po7119, po7120, po7121, po7122, po7123, po7124, po7125,
    po7126, po7127, po7128, po7129, po7130, po7131, po7132, po7133, po7134,
    po7135, po7136, po7137, po7138, po7139, po7140, po7141, po7142, po7143,
    po7144, po7145, po7146, po7147, po7148, po7149, po7150, po7151, po7152,
    po7153, po7154, po7155, po7156, po7157, po7158, po7159, po7160, po7161,
    po7162, po7163, po7164, po7165;
  wire new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294,
    new_n4295, new_n4296, new_n4297, new_n4298, new_n4299, new_n4300,
    new_n4301, new_n4302, new_n4303, new_n4304, new_n4305, new_n4306,
    new_n4307, new_n4308, new_n4309, new_n4310, new_n4311, new_n4312,
    new_n4313, new_n4314, new_n4315, new_n4316, new_n4317, new_n4318,
    new_n4319, new_n4320, new_n4321, new_n4322, new_n4323, new_n4324,
    new_n4325, new_n4326, new_n4327, new_n4328, new_n4329, new_n4330,
    new_n4331, new_n4332, new_n4333, new_n4334, new_n4335, new_n4336,
    new_n4337, new_n4338, new_n4339, new_n4340, new_n4341, new_n4342,
    new_n4343, new_n4344, new_n4345, new_n4346, new_n4347, new_n4348,
    new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354,
    new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360,
    new_n4361, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366,
    new_n4367, new_n4368, new_n4369, new_n4370, new_n4371, new_n4372,
    new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378,
    new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384,
    new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390,
    new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396,
    new_n4397, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402,
    new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408,
    new_n4409, new_n4410, new_n4411, new_n4412, new_n4413, new_n4414,
    new_n4415, new_n4416, new_n4417, new_n4418, new_n4419, new_n4420,
    new_n4421, new_n4422, new_n4423, new_n4424, new_n4425, new_n4426,
    new_n4427, new_n4428, new_n4429, new_n4430, new_n4431, new_n4432,
    new_n4433, new_n4434, new_n4435, new_n4436, new_n4437, new_n4438,
    new_n4439, new_n4440, new_n4441, new_n4442, new_n4443, new_n4444,
    new_n4445, new_n4446, new_n4447, new_n4448, new_n4449, new_n4450,
    new_n4451, new_n4452, new_n4453, new_n4454, new_n4455, new_n4456,
    new_n4457, new_n4458, new_n4459, new_n4460, new_n4461, new_n4462,
    new_n4463, new_n4464, new_n4465, new_n4466, new_n4467, new_n4468,
    new_n4469, new_n4470, new_n4471, new_n4472, new_n4473, new_n4474,
    new_n4475, new_n4476, new_n4477, new_n4478, new_n4479, new_n4480,
    new_n4481, new_n4482, new_n4483, new_n4484, new_n4485, new_n4486,
    new_n4487, new_n4488, new_n4489, new_n4490, new_n4491, new_n4492,
    new_n4493, new_n4494, new_n4495, new_n4496, new_n4497, new_n4498,
    new_n4499, new_n4500, new_n4501, new_n4502, new_n4503, new_n4504,
    new_n4505, new_n4506, new_n4507, new_n4508, new_n4509, new_n4510,
    new_n4511, new_n4512, new_n4513, new_n4514, new_n4515, new_n4516,
    new_n4517, new_n4518, new_n4519, new_n4520, new_n4521, new_n4522,
    new_n4523, new_n4524, new_n4525, new_n4526, new_n4527, new_n4528,
    new_n4529, new_n4530, new_n4531, new_n4532, new_n4533, new_n4534,
    new_n4535, new_n4536, new_n4537, new_n4538, new_n4539, new_n4540,
    new_n4541, new_n4542, new_n4543, new_n4544, new_n4545, new_n4546,
    new_n4547, new_n4548, new_n4549, new_n4550, new_n4551, new_n4552,
    new_n4553, new_n4554, new_n4555, new_n4556, new_n4557, new_n4558,
    new_n4559, new_n4560, new_n4561, new_n4562, new_n4563, new_n4564,
    new_n4565, new_n4566, new_n4567, new_n4568, new_n4569, new_n4570,
    new_n4571, new_n4572, new_n4573, new_n4574, new_n4575, new_n4576,
    new_n4577, new_n4578, new_n4579, new_n4580, new_n4581, new_n4582,
    new_n4583, new_n4584, new_n4585, new_n4586, new_n4587, new_n4588,
    new_n4589, new_n4590, new_n4591, new_n4592, new_n4593, new_n4594,
    new_n4595, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618,
    new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624,
    new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630,
    new_n4631, new_n4632, new_n4633, new_n4634, new_n4635, new_n4636,
    new_n4637, new_n4638, new_n4639, new_n4640, new_n4641, new_n4642,
    new_n4643, new_n4644, new_n4645, new_n4646, new_n4647, new_n4648,
    new_n4649, new_n4650, new_n4651, new_n4652, new_n4653, new_n4654,
    new_n4655, new_n4656, new_n4657, new_n4658, new_n4659, new_n4660,
    new_n4661, new_n4662, new_n4663, new_n4664, new_n4665, new_n4666,
    new_n4667, new_n4668, new_n4669, new_n4670, new_n4671, new_n4672,
    new_n4673, new_n4674, new_n4675, new_n4676, new_n4677, new_n4678,
    new_n4679, new_n4680, new_n4681, new_n4682, new_n4683, new_n4684,
    new_n4685, new_n4686, new_n4687, new_n4688, new_n4689, new_n4690,
    new_n4691, new_n4692, new_n4693, new_n4694, new_n4695, new_n4696,
    new_n4697, new_n4698, new_n4699, new_n4700, new_n4701, new_n4702,
    new_n4703, new_n4704, new_n4705, new_n4706, new_n4707, new_n4708,
    new_n4709, new_n4710, new_n4711, new_n4712, new_n4713, new_n4714,
    new_n4715, new_n4716, new_n4717, new_n4718, new_n4719, new_n4720,
    new_n4721, new_n4722, new_n4723, new_n4724, new_n4725, new_n4726,
    new_n4727, new_n4728, new_n4729, new_n4730, new_n4731, new_n4732,
    new_n4733, new_n4734, new_n4735, new_n4736, new_n4737, new_n4738,
    new_n4739, new_n4740, new_n4741, new_n4742, new_n4743, new_n4744,
    new_n4745, new_n4746, new_n4747, new_n4748, new_n4749, new_n4750,
    new_n4751, new_n4752, new_n4753, new_n4754, new_n4755, new_n4756,
    new_n4757, new_n4758, new_n4759, new_n4760, new_n4761, new_n4762,
    new_n4763, new_n4764, new_n4765, new_n4766, new_n4767, new_n4768,
    new_n4769, new_n4770, new_n4771, new_n4772, new_n4773, new_n4774,
    new_n4775, new_n4776, new_n4777, new_n4778, new_n4779, new_n4780,
    new_n4781, new_n4782, new_n4783, new_n4784, new_n4785, new_n4786,
    new_n4787, new_n4788, new_n4789, new_n4790, new_n4791, new_n4792,
    new_n4793, new_n4794, new_n4795, new_n4796, new_n4797, new_n4798,
    new_n4799, new_n4800, new_n4801, new_n4802, new_n4803, new_n4804,
    new_n4805, new_n4806, new_n4807, new_n4808, new_n4809, new_n4810,
    new_n4811, new_n4812, new_n4813, new_n4814, new_n4815, new_n4816,
    new_n4817, new_n4818, new_n4819, new_n4820, new_n4821, new_n4822,
    new_n4823, new_n4824, new_n4825, new_n4826, new_n4827, new_n4828,
    new_n4829, new_n4830, new_n4831, new_n4832, new_n4833, new_n4834,
    new_n4835, new_n4836, new_n4837, new_n4838, new_n4839, new_n4840,
    new_n4841, new_n4842, new_n4843, new_n4844, new_n4845, new_n4846,
    new_n4847, new_n4848, new_n4849, new_n4850, new_n4851, new_n4852,
    new_n4853, new_n4854, new_n4855, new_n4856, new_n4857, new_n4858,
    new_n4859, new_n4860, new_n4861, new_n4862, new_n4863, new_n4864,
    new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870,
    new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876,
    new_n4877, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882,
    new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888,
    new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894,
    new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948,
    new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954,
    new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960,
    new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966,
    new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972,
    new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978,
    new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990,
    new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996,
    new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644,
    new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693, new_n5694, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6005, new_n6006, new_n6007, new_n6008, new_n6009, new_n6010,
    new_n6011, new_n6012, new_n6013, new_n6014, new_n6015, new_n6016,
    new_n6017, new_n6018, new_n6019, new_n6020, new_n6021, new_n6022,
    new_n6023, new_n6024, new_n6025, new_n6026, new_n6027, new_n6028,
    new_n6029, new_n6030, new_n6031, new_n6032, new_n6033, new_n6034,
    new_n6035, new_n6036, new_n6037, new_n6038, new_n6039, new_n6040,
    new_n6041, new_n6042, new_n6043, new_n6044, new_n6045, new_n6046,
    new_n6047, new_n6048, new_n6049, new_n6050, new_n6051, new_n6052,
    new_n6053, new_n6054, new_n6055, new_n6056, new_n6057, new_n6058,
    new_n6059, new_n6060, new_n6061, new_n6062, new_n6063, new_n6064,
    new_n6065, new_n6066, new_n6067, new_n6068, new_n6069, new_n6070,
    new_n6071, new_n6072, new_n6073, new_n6074, new_n6075, new_n6076,
    new_n6077, new_n6078, new_n6079, new_n6080, new_n6081, new_n6082,
    new_n6083, new_n6084, new_n6085, new_n6086, new_n6087, new_n6088,
    new_n6089, new_n6090, new_n6091, new_n6092, new_n6093, new_n6094,
    new_n6095, new_n6096, new_n6097, new_n6098, new_n6099, new_n6100,
    new_n6101, new_n6102, new_n6103, new_n6104, new_n6105, new_n6106,
    new_n6107, new_n6108, new_n6109, new_n6110, new_n6111, new_n6112,
    new_n6113, new_n6114, new_n6115, new_n6116, new_n6117, new_n6118,
    new_n6119, new_n6120, new_n6121, new_n6122, new_n6123, new_n6124,
    new_n6125, new_n6126, new_n6127, new_n6128, new_n6129, new_n6130,
    new_n6131, new_n6132, new_n6133, new_n6134, new_n6135, new_n6136,
    new_n6137, new_n6138, new_n6139, new_n6140, new_n6141, new_n6142,
    new_n6143, new_n6144, new_n6145, new_n6146, new_n6147, new_n6148,
    new_n6149, new_n6150, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160,
    new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166,
    new_n6167, new_n6168, new_n6169, new_n6170, new_n6171, new_n6172,
    new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178,
    new_n6179, new_n6180, new_n6181, new_n6182, new_n6183, new_n6184,
    new_n6185, new_n6186, new_n6187, new_n6188, new_n6189, new_n6190,
    new_n6191, new_n6192, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204, new_n6205, new_n6206, new_n6207, new_n6208,
    new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214,
    new_n6215, new_n6216, new_n6217, new_n6218, new_n6219, new_n6220,
    new_n6221, new_n6222, new_n6223, new_n6224, new_n6225, new_n6226,
    new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232,
    new_n6233, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238,
    new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6244,
    new_n6245, new_n6246, new_n6247, new_n6248, new_n6249, new_n6250,
    new_n6251, new_n6252, new_n6253, new_n6254, new_n6255, new_n6256,
    new_n6257, new_n6258, new_n6259, new_n6260, new_n6261, new_n6262,
    new_n6263, new_n6264, new_n6265, new_n6266, new_n6267, new_n6268,
    new_n6269, new_n6270, new_n6271, new_n6272, new_n6273, new_n6274,
    new_n6275, new_n6276, new_n6277, new_n6278, new_n6279, new_n6280,
    new_n6281, new_n6282, new_n6283, new_n6284, new_n6285, new_n6286,
    new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292,
    new_n6293, new_n6294, new_n6295, new_n6296, new_n6297, new_n6298,
    new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304,
    new_n6305, new_n6306, new_n6307, new_n6308, new_n6309, new_n6310,
    new_n6311, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316,
    new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322,
    new_n6323, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328,
    new_n6329, new_n6330, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354, new_n6355, new_n6356, new_n6357, new_n6358,
    new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375, new_n6376,
    new_n6377, new_n6378, new_n6379, new_n6380, new_n6381, new_n6382,
    new_n6383, new_n6384, new_n6385, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427, new_n6428, new_n6429, new_n6430,
    new_n6431, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442,
    new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472,
    new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478,
    new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502,
    new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514,
    new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542, new_n6543, new_n6544,
    new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550,
    new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556,
    new_n6557, new_n6558, new_n6559, new_n6560, new_n6561, new_n6562,
    new_n6563, new_n6564, new_n6565, new_n6566, new_n6567, new_n6568,
    new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574,
    new_n6575, new_n6576, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586,
    new_n6587, new_n6588, new_n6589, new_n6590, new_n6591, new_n6592,
    new_n6593, new_n6594, new_n6595, new_n6596, new_n6597, new_n6598,
    new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604,
    new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6610,
    new_n6611, new_n6612, new_n6613, new_n6614, new_n6615, new_n6616,
    new_n6617, new_n6618, new_n6619, new_n6620, new_n6621, new_n6622,
    new_n6623, new_n6624, new_n6625, new_n6626, new_n6627, new_n6628,
    new_n6629, new_n6630, new_n6631, new_n6632, new_n6633, new_n6634,
    new_n6635, new_n6636, new_n6637, new_n6638, new_n6639, new_n6640,
    new_n6641, new_n6642, new_n6643, new_n6644, new_n6645, new_n6646,
    new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652,
    new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658,
    new_n6659, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664,
    new_n6665, new_n6666, new_n6667, new_n6668, new_n6669, new_n6670,
    new_n6671, new_n6672, new_n6673, new_n6674, new_n6675, new_n6676,
    new_n6677, new_n6678, new_n6679, new_n6680, new_n6681, new_n6682,
    new_n6683, new_n6684, new_n6685, new_n6686, new_n6687, new_n6688,
    new_n6689, new_n6690, new_n6691, new_n6692, new_n6693, new_n6694,
    new_n6695, new_n6696, new_n6697, new_n6698, new_n6699, new_n6700,
    new_n6701, new_n6702, new_n6703, new_n6704, new_n6705, new_n6706,
    new_n6707, new_n6708, new_n6709, new_n6710, new_n6711, new_n6712,
    new_n6713, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718,
    new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724,
    new_n6725, new_n6726, new_n6727, new_n6728, new_n6729, new_n6730,
    new_n6731, new_n6732, new_n6733, new_n6734, new_n6735, new_n6736,
    new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742,
    new_n6743, new_n6744, new_n6745, new_n6746, new_n6747, new_n6748,
    new_n6749, new_n6750, new_n6751, new_n6752, new_n6753, new_n6754,
    new_n6755, new_n6756, new_n6757, new_n6758, new_n6759, new_n6760,
    new_n6761, new_n6762, new_n6763, new_n6764, new_n6765, new_n6766,
    new_n6767, new_n6768, new_n6769, new_n6770, new_n6771, new_n6772,
    new_n6773, new_n6774, new_n6775, new_n6776, new_n6777, new_n6778,
    new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784,
    new_n6785, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790,
    new_n6791, new_n6792, new_n6793, new_n6794, new_n6795, new_n6796,
    new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802,
    new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808,
    new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814,
    new_n6815, new_n6816, new_n6817, new_n6818, new_n6819, new_n6820,
    new_n6821, new_n6822, new_n6823, new_n6824, new_n6825, new_n6826,
    new_n6827, new_n6828, new_n6829, new_n6830, new_n6831, new_n6832,
    new_n6833, new_n6834, new_n6835, new_n6836, new_n6837, new_n6838,
    new_n6839, new_n6840, new_n6841, new_n6842, new_n6843, new_n6844,
    new_n6845, new_n6846, new_n6847, new_n6848, new_n6849, new_n6850,
    new_n6851, new_n6852, new_n6853, new_n6854, new_n6855, new_n6856,
    new_n6857, new_n6858, new_n6859, new_n6860, new_n6861, new_n6862,
    new_n6863, new_n6864, new_n6865, new_n6866, new_n6867, new_n6868,
    new_n6869, new_n6870, new_n6871, new_n6872, new_n6873, new_n6874,
    new_n6875, new_n6876, new_n6877, new_n6878, new_n6879, new_n6880,
    new_n6881, new_n6882, new_n6883, new_n6884, new_n6885, new_n6886,
    new_n6887, new_n6888, new_n6889, new_n6890, new_n6891, new_n6892,
    new_n6893, new_n6894, new_n6895, new_n6896, new_n6897, new_n6898,
    new_n6899, new_n6900, new_n6901, new_n6902, new_n6903, new_n6904,
    new_n6905, new_n6906, new_n6907, new_n6908, new_n6909, new_n6910,
    new_n6911, new_n6912, new_n6913, new_n6914, new_n6915, new_n6916,
    new_n6917, new_n6918, new_n6919, new_n6920, new_n6921, new_n6922,
    new_n6923, new_n6924, new_n6925, new_n6926, new_n6927, new_n6928,
    new_n6929, new_n6930, new_n6931, new_n6932, new_n6933, new_n6934,
    new_n6935, new_n6936, new_n6937, new_n6938, new_n6939, new_n6940,
    new_n6941, new_n6942, new_n6943, new_n6944, new_n6945, new_n6946,
    new_n6947, new_n6948, new_n6949, new_n6950, new_n6951, new_n6952,
    new_n6953, new_n6954, new_n6955, new_n6956, new_n6957, new_n6958,
    new_n6959, new_n6960, new_n6961, new_n6962, new_n6963, new_n6964,
    new_n6965, new_n6966, new_n6967, new_n6968, new_n6969, new_n6970,
    new_n6971, new_n6972, new_n6973, new_n6974, new_n6975, new_n6976,
    new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982,
    new_n6983, new_n6984, new_n6985, new_n6986, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072,
    new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078,
    new_n7079, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084,
    new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090,
    new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096,
    new_n7097, new_n7098, new_n7099, new_n7100, new_n7101, new_n7102,
    new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108,
    new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114,
    new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120,
    new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190, new_n7191, new_n7192,
    new_n7193, new_n7194, new_n7195, new_n7196, new_n7197, new_n7198,
    new_n7199, new_n7200, new_n7201, new_n7202, new_n7203, new_n7204,
    new_n7205, new_n7206, new_n7207, new_n7208, new_n7209, new_n7210,
    new_n7211, new_n7212, new_n7213, new_n7214, new_n7215, new_n7216,
    new_n7217, new_n7218, new_n7219, new_n7220, new_n7221, new_n7222,
    new_n7223, new_n7224, new_n7225, new_n7226, new_n7227, new_n7228,
    new_n7229, new_n7230, new_n7231, new_n7232, new_n7233, new_n7234,
    new_n7235, new_n7236, new_n7237, new_n7238, new_n7239, new_n7240,
    new_n7241, new_n7242, new_n7243, new_n7244, new_n7245, new_n7246,
    new_n7247, new_n7248, new_n7249, new_n7250, new_n7251, new_n7252,
    new_n7253, new_n7254, new_n7255, new_n7256, new_n7257, new_n7258,
    new_n7259, new_n7260, new_n7261, new_n7262, new_n7263, new_n7264,
    new_n7265, new_n7266, new_n7267, new_n7268, new_n7269, new_n7270,
    new_n7271, new_n7272, new_n7273, new_n7274, new_n7275, new_n7276,
    new_n7277, new_n7278, new_n7279, new_n7280, new_n7281, new_n7282,
    new_n7283, new_n7284, new_n7285, new_n7286, new_n7287, new_n7288,
    new_n7289, new_n7290, new_n7291, new_n7292, new_n7293, new_n7294,
    new_n7295, new_n7296, new_n7297, new_n7298, new_n7299, new_n7300,
    new_n7301, new_n7302, new_n7303, new_n7304, new_n7305, new_n7306,
    new_n7307, new_n7308, new_n7309, new_n7310, new_n7311, new_n7312,
    new_n7313, new_n7314, new_n7315, new_n7316, new_n7317, new_n7318,
    new_n7319, new_n7320, new_n7321, new_n7322, new_n7323, new_n7324,
    new_n7325, new_n7326, new_n7327, new_n7328, new_n7329, new_n7330,
    new_n7331, new_n7332, new_n7333, new_n7334, new_n7335, new_n7336,
    new_n7337, new_n7338, new_n7339, new_n7340, new_n7341, new_n7342,
    new_n7343, new_n7344, new_n7345, new_n7346, new_n7347, new_n7348,
    new_n7349, new_n7350, new_n7351, new_n7352, new_n7353, new_n7354,
    new_n7355, new_n7356, new_n7357, new_n7358, new_n7359, new_n7360,
    new_n7361, new_n7362, new_n7363, new_n7364, new_n7365, new_n7366,
    new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372,
    new_n7373, new_n7374, new_n7375, new_n7376, new_n7377, new_n7378,
    new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384,
    new_n7385, new_n7386, new_n7387, new_n7388, new_n7389, new_n7390,
    new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396,
    new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402,
    new_n7403, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408,
    new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7414,
    new_n7415, new_n7416, new_n7417, new_n7418, new_n7419, new_n7420,
    new_n7421, new_n7422, new_n7423, new_n7424, new_n7425, new_n7426,
    new_n7427, new_n7428, new_n7429, new_n7430, new_n7431, new_n7432,
    new_n7433, new_n7434, new_n7435, new_n7436, new_n7437, new_n7438,
    new_n7439, new_n7440, new_n7441, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456,
    new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566, new_n7567, new_n7568, new_n7569, new_n7570,
    new_n7571, new_n7572, new_n7573, new_n7574, new_n7575, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585, new_n7586, new_n7587, new_n7588,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607, new_n7608, new_n7609, new_n7610, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616, new_n7617, new_n7618,
    new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624,
    new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630,
    new_n7631, new_n7632, new_n7633, new_n7634, new_n7635, new_n7636,
    new_n7637, new_n7638, new_n7639, new_n7640, new_n7641, new_n7642,
    new_n7643, new_n7644, new_n7645, new_n7646, new_n7647, new_n7648,
    new_n7649, new_n7650, new_n7651, new_n7652, new_n7653, new_n7654,
    new_n7655, new_n7656, new_n7657, new_n7658, new_n7659, new_n7660,
    new_n7661, new_n7662, new_n7663, new_n7664, new_n7665, new_n7666,
    new_n7667, new_n7668, new_n7669, new_n7670, new_n7671, new_n7672,
    new_n7673, new_n7674, new_n7675, new_n7676, new_n7677, new_n7678,
    new_n7679, new_n7680, new_n7681, new_n7682, new_n7683, new_n7684,
    new_n7685, new_n7686, new_n7687, new_n7688, new_n7689, new_n7690,
    new_n7691, new_n7692, new_n7693, new_n7694, new_n7695, new_n7696,
    new_n7697, new_n7698, new_n7699, new_n7700, new_n7701, new_n7702,
    new_n7703, new_n7704, new_n7705, new_n7706, new_n7707, new_n7708,
    new_n7709, new_n7710, new_n7711, new_n7712, new_n7713, new_n7714,
    new_n7715, new_n7716, new_n7717, new_n7718, new_n7719, new_n7720,
    new_n7721, new_n7722, new_n7723, new_n7724, new_n7725, new_n7726,
    new_n7727, new_n7728, new_n7729, new_n7730, new_n7731, new_n7732,
    new_n7733, new_n7734, new_n7735, new_n7736, new_n7737, new_n7738,
    new_n7739, new_n7740, new_n7741, new_n7742, new_n7743, new_n7744,
    new_n7745, new_n7746, new_n7747, new_n7748, new_n7749, new_n7750,
    new_n7751, new_n7752, new_n7753, new_n7754, new_n7755, new_n7756,
    new_n7757, new_n7758, new_n7759, new_n7760, new_n7761, new_n7762,
    new_n7763, new_n7764, new_n7765, new_n7766, new_n7767, new_n7768,
    new_n7769, new_n7770, new_n7771, new_n7772, new_n7773, new_n7774,
    new_n7775, new_n7776, new_n7777, new_n7778, new_n7779, new_n7780,
    new_n7781, new_n7782, new_n7783, new_n7784, new_n7785, new_n7786,
    new_n7787, new_n7788, new_n7789, new_n7790, new_n7791, new_n7792,
    new_n7793, new_n7794, new_n7795, new_n7796, new_n7797, new_n7798,
    new_n7799, new_n7800, new_n7801, new_n7802, new_n7803, new_n7804,
    new_n7805, new_n7806, new_n7807, new_n7808, new_n7809, new_n7810,
    new_n7811, new_n7812, new_n7813, new_n7814, new_n7815, new_n7816,
    new_n7817, new_n7818, new_n7819, new_n7820, new_n7821, new_n7822,
    new_n7823, new_n7824, new_n7825, new_n7826, new_n7827, new_n7828,
    new_n7829, new_n7830, new_n7831, new_n7832, new_n7833, new_n7834,
    new_n7835, new_n7836, new_n7837, new_n7838, new_n7839, new_n7840,
    new_n7841, new_n7842, new_n7843, new_n7844, new_n7845, new_n7846,
    new_n7847, new_n7848, new_n7849, new_n7850, new_n7851, new_n7852,
    new_n7853, new_n7854, new_n7855, new_n7856, new_n7857, new_n7858,
    new_n7859, new_n7860, new_n7861, new_n7862, new_n7863, new_n7864,
    new_n7865, new_n7866, new_n7867, new_n7868, new_n7869, new_n7870,
    new_n7871, new_n7872, new_n7873, new_n7874, new_n7875, new_n7876,
    new_n7877, new_n7878, new_n7879, new_n7880, new_n7881, new_n7882,
    new_n7883, new_n7884, new_n7885, new_n7886, new_n7887, new_n7888,
    new_n7889, new_n7890, new_n7891, new_n7892, new_n7893, new_n7894,
    new_n7895, new_n7896, new_n7897, new_n7898, new_n7899, new_n7900,
    new_n7901, new_n7902, new_n7903, new_n7904, new_n7905, new_n7906,
    new_n7907, new_n7908, new_n7909, new_n7910, new_n7911, new_n7912,
    new_n7913, new_n7914, new_n7915, new_n7916, new_n7917, new_n7918,
    new_n7919, new_n7920, new_n7921, new_n7922, new_n7923, new_n7924,
    new_n7925, new_n7926, new_n7927, new_n7928, new_n7929, new_n7930,
    new_n7931, new_n7932, new_n7933, new_n7934, new_n7935, new_n7936,
    new_n7937, new_n7938, new_n7939, new_n7940, new_n7941, new_n7942,
    new_n7943, new_n7944, new_n7945, new_n7946, new_n7947, new_n7948,
    new_n7949, new_n7950, new_n7951, new_n7952, new_n7953, new_n7954,
    new_n7955, new_n7956, new_n7957, new_n7958, new_n7959, new_n7960,
    new_n7961, new_n7962, new_n7963, new_n7964, new_n7965, new_n7966,
    new_n7967, new_n7968, new_n7969, new_n7970, new_n7971, new_n7972,
    new_n7973, new_n7974, new_n7975, new_n7976, new_n7977, new_n7978,
    new_n7979, new_n7980, new_n7981, new_n7982, new_n7983, new_n7984,
    new_n7985, new_n7986, new_n7987, new_n7988, new_n7989, new_n7990,
    new_n7991, new_n7992, new_n7993, new_n7994, new_n7995, new_n7996,
    new_n7997, new_n7998, new_n7999, new_n8000, new_n8001, new_n8002,
    new_n8003, new_n8004, new_n8005, new_n8006, new_n8007, new_n8008,
    new_n8009, new_n8010, new_n8011, new_n8012, new_n8013, new_n8014,
    new_n8015, new_n8016, new_n8017, new_n8018, new_n8019, new_n8020,
    new_n8021, new_n8022, new_n8023, new_n8024, new_n8025, new_n8026,
    new_n8027, new_n8028, new_n8029, new_n8030, new_n8031, new_n8032,
    new_n8033, new_n8034, new_n8035, new_n8036, new_n8037, new_n8038,
    new_n8039, new_n8040, new_n8041, new_n8042, new_n8043, new_n8044,
    new_n8045, new_n8046, new_n8047, new_n8048, new_n8049, new_n8050,
    new_n8051, new_n8052, new_n8053, new_n8054, new_n8055, new_n8056,
    new_n8057, new_n8058, new_n8059, new_n8060, new_n8061, new_n8062,
    new_n8063, new_n8064, new_n8065, new_n8066, new_n8067, new_n8068,
    new_n8069, new_n8070, new_n8071, new_n8072, new_n8073, new_n8074,
    new_n8075, new_n8076, new_n8077, new_n8078, new_n8079, new_n8080,
    new_n8081, new_n8082, new_n8083, new_n8084, new_n8085, new_n8086,
    new_n8087, new_n8088, new_n8089, new_n8090, new_n8091, new_n8092,
    new_n8093, new_n8094, new_n8095, new_n8096, new_n8097, new_n8098,
    new_n8099, new_n8100, new_n8101, new_n8102, new_n8103, new_n8104,
    new_n8105, new_n8106, new_n8107, new_n8108, new_n8109, new_n8110,
    new_n8111, new_n8112, new_n8113, new_n8114, new_n8115, new_n8116,
    new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122,
    new_n8123, new_n8124, new_n8125, new_n8126, new_n8127, new_n8128,
    new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134,
    new_n8135, new_n8136, new_n8137, new_n8138, new_n8139, new_n8140,
    new_n8141, new_n8142, new_n8143, new_n8144, new_n8145, new_n8146,
    new_n8147, new_n8148, new_n8149, new_n8150, new_n8151, new_n8152,
    new_n8153, new_n8154, new_n8155, new_n8156, new_n8157, new_n8158,
    new_n8159, new_n8160, new_n8161, new_n8162, new_n8163, new_n8164,
    new_n8165, new_n8166, new_n8167, new_n8168, new_n8169, new_n8170,
    new_n8171, new_n8172, new_n8173, new_n8174, new_n8175, new_n8176,
    new_n8177, new_n8178, new_n8179, new_n8180, new_n8181, new_n8182,
    new_n8183, new_n8184, new_n8185, new_n8186, new_n8187, new_n8188,
    new_n8189, new_n8190, new_n8191, new_n8192, new_n8193, new_n8194,
    new_n8195, new_n8196, new_n8197, new_n8198, new_n8199, new_n8200,
    new_n8201, new_n8202, new_n8203, new_n8204, new_n8205, new_n8206,
    new_n8207, new_n8208, new_n8209, new_n8210, new_n8211, new_n8212,
    new_n8213, new_n8214, new_n8215, new_n8216, new_n8217, new_n8218,
    new_n8219, new_n8220, new_n8221, new_n8222, new_n8223, new_n8224,
    new_n8225, new_n8226, new_n8227, new_n8228, new_n8229, new_n8230,
    new_n8231, new_n8232, new_n8233, new_n8234, new_n8235, new_n8236,
    new_n8237, new_n8238, new_n8239, new_n8240, new_n8241, new_n8242,
    new_n8243, new_n8244, new_n8245, new_n8246, new_n8247, new_n8248,
    new_n8249, new_n8250, new_n8251, new_n8252, new_n8253, new_n8254,
    new_n8255, new_n8256, new_n8257, new_n8258, new_n8259, new_n8260,
    new_n8261, new_n8262, new_n8263, new_n8264, new_n8265, new_n8266,
    new_n8267, new_n8268, new_n8269, new_n8270, new_n8271, new_n8272,
    new_n8273, new_n8274, new_n8275, new_n8276, new_n8277, new_n8278,
    new_n8279, new_n8280, new_n8281, new_n8282, new_n8283, new_n8284,
    new_n8285, new_n8286, new_n8287, new_n8288, new_n8289, new_n8290,
    new_n8291, new_n8292, new_n8293, new_n8294, new_n8295, new_n8296,
    new_n8297, new_n8298, new_n8299, new_n8300, new_n8301, new_n8302,
    new_n8303, new_n8304, new_n8305, new_n8306, new_n8307, new_n8308,
    new_n8309, new_n8310, new_n8311, new_n8312, new_n8313, new_n8314,
    new_n8315, new_n8316, new_n8317, new_n8318, new_n8319, new_n8320,
    new_n8321, new_n8322, new_n8323, new_n8324, new_n8325, new_n8326,
    new_n8327, new_n8328, new_n8329, new_n8330, new_n8331, new_n8332,
    new_n8333, new_n8334, new_n8335, new_n8336, new_n8337, new_n8338,
    new_n8339, new_n8340, new_n8341, new_n8342, new_n8343, new_n8344,
    new_n8345, new_n8346, new_n8347, new_n8348, new_n8349, new_n8350,
    new_n8351, new_n8352, new_n8353, new_n8354, new_n8355, new_n8356,
    new_n8357, new_n8358, new_n8359, new_n8360, new_n8361, new_n8362,
    new_n8363, new_n8364, new_n8365, new_n8366, new_n8367, new_n8368,
    new_n8369, new_n8370, new_n8371, new_n8372, new_n8373, new_n8374,
    new_n8375, new_n8376, new_n8377, new_n8378, new_n8379, new_n8380,
    new_n8381, new_n8382, new_n8383, new_n8384, new_n8385, new_n8386,
    new_n8387, new_n8388, new_n8389, new_n8390, new_n8391, new_n8392,
    new_n8393, new_n8394, new_n8395, new_n8396, new_n8397, new_n8398,
    new_n8399, new_n8400, new_n8401, new_n8402, new_n8403, new_n8404,
    new_n8405, new_n8406, new_n8407, new_n8408, new_n8409, new_n8410,
    new_n8411, new_n8412, new_n8413, new_n8414, new_n8415, new_n8416,
    new_n8417, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422,
    new_n8423, new_n8424, new_n8425, new_n8426, new_n8427, new_n8428,
    new_n8429, new_n8430, new_n8431, new_n8432, new_n8433, new_n8434,
    new_n8435, new_n8436, new_n8437, new_n8438, new_n8439, new_n8440,
    new_n8441, new_n8442, new_n8443, new_n8444, new_n8445, new_n8446,
    new_n8447, new_n8448, new_n8449, new_n8450, new_n8451, new_n8452,
    new_n8453, new_n8454, new_n8455, new_n8456, new_n8457, new_n8458,
    new_n8459, new_n8460, new_n8461, new_n8462, new_n8463, new_n8464,
    new_n8465, new_n8466, new_n8467, new_n8468, new_n8469, new_n8470,
    new_n8471, new_n8472, new_n8473, new_n8474, new_n8475, new_n8476,
    new_n8477, new_n8478, new_n8479, new_n8480, new_n8481, new_n8482,
    new_n8483, new_n8484, new_n8485, new_n8486, new_n8487, new_n8488,
    new_n8489, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494,
    new_n8495, new_n8496, new_n8497, new_n8498, new_n8499, new_n8500,
    new_n8501, new_n8502, new_n8503, new_n8504, new_n8505, new_n8506,
    new_n8507, new_n8508, new_n8509, new_n8510, new_n8511, new_n8512,
    new_n8513, new_n8514, new_n8515, new_n8516, new_n8517, new_n8518,
    new_n8519, new_n8520, new_n8521, new_n8522, new_n8523, new_n8524,
    new_n8525, new_n8526, new_n8527, new_n8528, new_n8529, new_n8530,
    new_n8531, new_n8532, new_n8533, new_n8534, new_n8535, new_n8536,
    new_n8537, new_n8538, new_n8539, new_n8540, new_n8541, new_n8542,
    new_n8543, new_n8544, new_n8545, new_n8546, new_n8547, new_n8548,
    new_n8549, new_n8550, new_n8551, new_n8552, new_n8553, new_n8554,
    new_n8555, new_n8556, new_n8557, new_n8558, new_n8559, new_n8560,
    new_n8561, new_n8562, new_n8563, new_n8564, new_n8565, new_n8566,
    new_n8567, new_n8568, new_n8569, new_n8570, new_n8571, new_n8572,
    new_n8573, new_n8574, new_n8575, new_n8576, new_n8577, new_n8578,
    new_n8579, new_n8580, new_n8581, new_n8582, new_n8583, new_n8584,
    new_n8585, new_n8586, new_n8587, new_n8588, new_n8589, new_n8590,
    new_n8591, new_n8592, new_n8593, new_n8594, new_n8595, new_n8596,
    new_n8597, new_n8598, new_n8599, new_n8600, new_n8601, new_n8602,
    new_n8603, new_n8604, new_n8605, new_n8606, new_n8607, new_n8608,
    new_n8609, new_n8610, new_n8611, new_n8612, new_n8613, new_n8614,
    new_n8615, new_n8616, new_n8617, new_n8618, new_n8619, new_n8620,
    new_n8621, new_n8622, new_n8623, new_n8624, new_n8625, new_n8626,
    new_n8627, new_n8628, new_n8629, new_n8630, new_n8631, new_n8632,
    new_n8633, new_n8634, new_n8635, new_n8636, new_n8637, new_n8638,
    new_n8639, new_n8640, new_n8641, new_n8642, new_n8643, new_n8644,
    new_n8645, new_n8646, new_n8647, new_n8648, new_n8649, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662,
    new_n8663, new_n8664, new_n8665, new_n8666, new_n8667, new_n8668,
    new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674,
    new_n8675, new_n8676, new_n8677, new_n8678, new_n8679, new_n8680,
    new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686,
    new_n8687, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692,
    new_n8693, new_n8694, new_n8695, new_n8696, new_n8697, new_n8698,
    new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704,
    new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710,
    new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716,
    new_n8717, new_n8718, new_n8719, new_n8720, new_n8721, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744, new_n8745, new_n8746,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803, new_n8804, new_n8805, new_n8806,
    new_n8807, new_n8808, new_n8809, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819, new_n8820, new_n8821, new_n8822, new_n8823, new_n8824,
    new_n8825, new_n8826, new_n8827, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861, new_n8862, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884,
    new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890,
    new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896,
    new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902,
    new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908,
    new_n8909, new_n8910, new_n8911, new_n8912, new_n8913, new_n8914,
    new_n8915, new_n8916, new_n8917, new_n8918, new_n8919, new_n8920,
    new_n8921, new_n8922, new_n8923, new_n8924, new_n8925, new_n8926,
    new_n8927, new_n8928, new_n8929, new_n8930, new_n8931, new_n8932,
    new_n8933, new_n8934, new_n8935, new_n8936, new_n8937, new_n8938,
    new_n8939, new_n8940, new_n8941, new_n8942, new_n8943, new_n8944,
    new_n8945, new_n8946, new_n8947, new_n8948, new_n8949, new_n8950,
    new_n8951, new_n8952, new_n8953, new_n8954, new_n8955, new_n8956,
    new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962,
    new_n8963, new_n8964, new_n8965, new_n8966, new_n8967, new_n8968,
    new_n8969, new_n8970, new_n8971, new_n8972, new_n8973, new_n8974,
    new_n8975, new_n8976, new_n8977, new_n8978, new_n8979, new_n8980,
    new_n8981, new_n8982, new_n8983, new_n8984, new_n8985, new_n8986,
    new_n8987, new_n8988, new_n8989, new_n8990, new_n8991, new_n8992,
    new_n8993, new_n8994, new_n8995, new_n8996, new_n8997, new_n8998,
    new_n8999, new_n9000, new_n9001, new_n9002, new_n9003, new_n9004,
    new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010,
    new_n9011, new_n9012, new_n9013, new_n9014, new_n9015, new_n9016,
    new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022,
    new_n9023, new_n9024, new_n9025, new_n9026, new_n9027, new_n9028,
    new_n9029, new_n9030, new_n9031, new_n9032, new_n9033, new_n9034,
    new_n9035, new_n9036, new_n9037, new_n9038, new_n9039, new_n9040,
    new_n9041, new_n9042, new_n9043, new_n9044, new_n9045, new_n9046,
    new_n9047, new_n9048, new_n9049, new_n9050, new_n9051, new_n9052,
    new_n9053, new_n9054, new_n9055, new_n9056, new_n9057, new_n9058,
    new_n9059, new_n9060, new_n9061, new_n9062, new_n9063, new_n9064,
    new_n9065, new_n9066, new_n9067, new_n9068, new_n9069, new_n9070,
    new_n9071, new_n9072, new_n9073, new_n9074, new_n9075, new_n9076,
    new_n9077, new_n9078, new_n9079, new_n9080, new_n9081, new_n9082,
    new_n9083, new_n9084, new_n9085, new_n9086, new_n9087, new_n9088,
    new_n9089, new_n9090, new_n9091, new_n9092, new_n9093, new_n9094,
    new_n9095, new_n9096, new_n9097, new_n9098, new_n9099, new_n9100,
    new_n9101, new_n9102, new_n9103, new_n9104, new_n9105, new_n9106,
    new_n9107, new_n9108, new_n9109, new_n9110, new_n9111, new_n9112,
    new_n9113, new_n9114, new_n9115, new_n9116, new_n9117, new_n9118,
    new_n9119, new_n9120, new_n9121, new_n9122, new_n9123, new_n9124,
    new_n9125, new_n9126, new_n9127, new_n9128, new_n9129, new_n9130,
    new_n9131, new_n9132, new_n9133, new_n9134, new_n9135, new_n9136,
    new_n9137, new_n9138, new_n9139, new_n9140, new_n9141, new_n9142,
    new_n9143, new_n9144, new_n9145, new_n9146, new_n9147, new_n9148,
    new_n9149, new_n9150, new_n9151, new_n9152, new_n9153, new_n9154,
    new_n9155, new_n9156, new_n9157, new_n9158, new_n9159, new_n9160,
    new_n9161, new_n9162, new_n9163, new_n9164, new_n9165, new_n9166,
    new_n9167, new_n9168, new_n9169, new_n9170, new_n9171, new_n9172,
    new_n9173, new_n9174, new_n9175, new_n9176, new_n9177, new_n9178,
    new_n9179, new_n9180, new_n9181, new_n9182, new_n9183, new_n9184,
    new_n9185, new_n9186, new_n9187, new_n9188, new_n9189, new_n9190,
    new_n9191, new_n9192, new_n9193, new_n9194, new_n9195, new_n9196,
    new_n9197, new_n9198, new_n9199, new_n9200, new_n9201, new_n9202,
    new_n9203, new_n9204, new_n9205, new_n9206, new_n9207, new_n9208,
    new_n9209, new_n9210, new_n9211, new_n9212, new_n9213, new_n9214,
    new_n9215, new_n9216, new_n9217, new_n9218, new_n9219, new_n9220,
    new_n9221, new_n9222, new_n9223, new_n9224, new_n9225, new_n9226,
    new_n9227, new_n9228, new_n9229, new_n9230, new_n9231, new_n9232,
    new_n9233, new_n9234, new_n9235, new_n9236, new_n9237, new_n9238,
    new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244,
    new_n9245, new_n9246, new_n9247, new_n9248, new_n9249, new_n9250,
    new_n9251, new_n9252, new_n9253, new_n9254, new_n9255, new_n9256,
    new_n9257, new_n9258, new_n9259, new_n9260, new_n9261, new_n9262,
    new_n9263, new_n9264, new_n9265, new_n9266, new_n9267, new_n9268,
    new_n9269, new_n9270, new_n9271, new_n9272, new_n9273, new_n9274,
    new_n9275, new_n9276, new_n9277, new_n9278, new_n9279, new_n9280,
    new_n9281, new_n9282, new_n9283, new_n9284, new_n9285, new_n9286,
    new_n9287, new_n9288, new_n9289, new_n9290, new_n9291, new_n9292,
    new_n9293, new_n9294, new_n9295, new_n9296, new_n9297, new_n9298,
    new_n9299, new_n9300, new_n9301, new_n9302, new_n9303, new_n9304,
    new_n9305, new_n9306, new_n9307, new_n9308, new_n9309, new_n9310,
    new_n9311, new_n9312, new_n9313, new_n9314, new_n9315, new_n9316,
    new_n9317, new_n9318, new_n9319, new_n9320, new_n9321, new_n9322,
    new_n9323, new_n9324, new_n9325, new_n9326, new_n9327, new_n9328,
    new_n9329, new_n9330, new_n9331, new_n9332, new_n9333, new_n9334,
    new_n9335, new_n9336, new_n9337, new_n9338, new_n9339, new_n9340,
    new_n9341, new_n9342, new_n9343, new_n9344, new_n9345, new_n9346,
    new_n9347, new_n9348, new_n9349, new_n9350, new_n9351, new_n9352,
    new_n9353, new_n9354, new_n9355, new_n9356, new_n9357, new_n9358,
    new_n9359, new_n9360, new_n9361, new_n9362, new_n9363, new_n9364,
    new_n9365, new_n9366, new_n9367, new_n9368, new_n9369, new_n9370,
    new_n9371, new_n9372, new_n9373, new_n9374, new_n9375, new_n9376,
    new_n9377, new_n9378, new_n9379, new_n9380, new_n9381, new_n9382,
    new_n9383, new_n9384, new_n9385, new_n9386, new_n9387, new_n9388,
    new_n9389, new_n9390, new_n9391, new_n9392, new_n9393, new_n9394,
    new_n9395, new_n9396, new_n9397, new_n9398, new_n9399, new_n9400,
    new_n9401, new_n9402, new_n9403, new_n9404, new_n9405, new_n9406,
    new_n9407, new_n9408, new_n9409, new_n9410, new_n9411, new_n9412,
    new_n9413, new_n9414, new_n9415, new_n9416, new_n9417, new_n9418,
    new_n9419, new_n9420, new_n9421, new_n9422, new_n9423, new_n9424,
    new_n9425, new_n9426, new_n9427, new_n9428, new_n9429, new_n9430,
    new_n9431, new_n9432, new_n9433, new_n9434, new_n9435, new_n9436,
    new_n9437, new_n9438, new_n9439, new_n9440, new_n9441, new_n9442,
    new_n9443, new_n9444, new_n9445, new_n9446, new_n9447, new_n9448,
    new_n9449, new_n9450, new_n9451, new_n9452, new_n9453, new_n9454,
    new_n9455, new_n9456, new_n9457, new_n9458, new_n9459, new_n9460,
    new_n9461, new_n9462, new_n9463, new_n9464, new_n9465, new_n9466,
    new_n9467, new_n9468, new_n9469, new_n9470, new_n9471, new_n9472,
    new_n9473, new_n9474, new_n9475, new_n9476, new_n9477, new_n9478,
    new_n9479, new_n9480, new_n9481, new_n9482, new_n9483, new_n9484,
    new_n9485, new_n9486, new_n9487, new_n9488, new_n9489, new_n9490,
    new_n9491, new_n9492, new_n9493, new_n9494, new_n9495, new_n9496,
    new_n9497, new_n9498, new_n9499, new_n9500, new_n9501, new_n9502,
    new_n9503, new_n9504, new_n9505, new_n9506, new_n9507, new_n9508,
    new_n9509, new_n9510, new_n9511, new_n9512, new_n9513, new_n9514,
    new_n9515, new_n9516, new_n9517, new_n9518, new_n9519, new_n9520,
    new_n9521, new_n9522, new_n9523, new_n9524, new_n9525, new_n9526,
    new_n9527, new_n9528, new_n9529, new_n9530, new_n9531, new_n9532,
    new_n9533, new_n9534, new_n9535, new_n9536, new_n9537, new_n9538,
    new_n9539, new_n9540, new_n9541, new_n9542, new_n9543, new_n9544,
    new_n9545, new_n9546, new_n9547, new_n9548, new_n9549, new_n9550,
    new_n9551, new_n9552, new_n9553, new_n9554, new_n9555, new_n9556,
    new_n9557, new_n9558, new_n9559, new_n9560, new_n9561, new_n9562,
    new_n9563, new_n9564, new_n9565, new_n9566, new_n9567, new_n9568,
    new_n9569, new_n9570, new_n9571, new_n9572, new_n9573, new_n9574,
    new_n9575, new_n9576, new_n9577, new_n9578, new_n9579, new_n9580,
    new_n9581, new_n9582, new_n9583, new_n9584, new_n9585, new_n9586,
    new_n9587, new_n9588, new_n9589, new_n9590, new_n9591, new_n9592,
    new_n9593, new_n9594, new_n9595, new_n9596, new_n9597, new_n9598,
    new_n9599, new_n9600, new_n9601, new_n9602, new_n9603, new_n9604,
    new_n9605, new_n9606, new_n9607, new_n9608, new_n9609, new_n9610,
    new_n9611, new_n9612, new_n9613, new_n9614, new_n9615, new_n9616,
    new_n9617, new_n9618, new_n9619, new_n9620, new_n9621, new_n9622,
    new_n9623, new_n9624, new_n9625, new_n9626, new_n9627, new_n9628,
    new_n9629, new_n9630, new_n9631, new_n9632, new_n9633, new_n9634,
    new_n9635, new_n9636, new_n9637, new_n9638, new_n9639, new_n9640,
    new_n9641, new_n9642, new_n9643, new_n9644, new_n9645, new_n9646,
    new_n9647, new_n9648, new_n9649, new_n9650, new_n9651, new_n9652,
    new_n9653, new_n9654, new_n9655, new_n9656, new_n9657, new_n9658,
    new_n9659, new_n9660, new_n9661, new_n9662, new_n9663, new_n9664,
    new_n9665, new_n9666, new_n9667, new_n9668, new_n9669, new_n9670,
    new_n9671, new_n9672, new_n9673, new_n9674, new_n9675, new_n9676,
    new_n9677, new_n9678, new_n9679, new_n9680, new_n9681, new_n9682,
    new_n9683, new_n9684, new_n9685, new_n9686, new_n9687, new_n9688,
    new_n9689, new_n9690, new_n9691, new_n9692, new_n9693, new_n9694,
    new_n9695, new_n9696, new_n9697, new_n9698, new_n9699, new_n9700,
    new_n9701, new_n9702, new_n9703, new_n9704, new_n9705, new_n9706,
    new_n9707, new_n9708, new_n9709, new_n9710, new_n9711, new_n9712,
    new_n9713, new_n9714, new_n9715, new_n9716, new_n9717, new_n9718,
    new_n9719, new_n9720, new_n9721, new_n9722, new_n9723, new_n9724,
    new_n9725, new_n9726, new_n9727, new_n9728, new_n9729, new_n9730,
    new_n9731, new_n9732, new_n9733, new_n9734, new_n9735, new_n9736,
    new_n9737, new_n9738, new_n9739, new_n9740, new_n9741, new_n9742,
    new_n9743, new_n9744, new_n9745, new_n9746, new_n9747, new_n9748,
    new_n9749, new_n9750, new_n9751, new_n9752, new_n9753, new_n9754,
    new_n9755, new_n9756, new_n9757, new_n9758, new_n9759, new_n9760,
    new_n9761, new_n9762, new_n9763, new_n9764, new_n9765, new_n9766,
    new_n9767, new_n9768, new_n9769, new_n9770, new_n9771, new_n9772,
    new_n9773, new_n9774, new_n9775, new_n9776, new_n9777, new_n9778,
    new_n9779, new_n9780, new_n9781, new_n9782, new_n9783, new_n9784,
    new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790,
    new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796,
    new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802,
    new_n9803, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808,
    new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814,
    new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820,
    new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826,
    new_n9827, new_n9828, new_n9829, new_n9830, new_n9831, new_n9832,
    new_n9833, new_n9834, new_n9835, new_n9836, new_n9837, new_n9838,
    new_n9839, new_n9840, new_n9841, new_n9842, new_n9843, new_n9844,
    new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850,
    new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856,
    new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862,
    new_n9863, new_n9864, new_n9865, new_n9866, new_n9867, new_n9868,
    new_n9869, new_n9870, new_n9871, new_n9872, new_n9873, new_n9874,
    new_n9875, new_n9876, new_n9877, new_n9878, new_n9879, new_n9880,
    new_n9881, new_n9882, new_n9883, new_n9884, new_n9885, new_n9886,
    new_n9887, new_n9888, new_n9889, new_n9890, new_n9891, new_n9892,
    new_n9893, new_n9894, new_n9895, new_n9896, new_n9897, new_n9898,
    new_n9899, new_n9900, new_n9901, new_n9902, new_n9903, new_n9904,
    new_n9905, new_n9906, new_n9907, new_n9908, new_n9909, new_n9910,
    new_n9911, new_n9912, new_n9913, new_n9914, new_n9915, new_n9916,
    new_n9917, new_n9918, new_n9919, new_n9920, new_n9921, new_n9922,
    new_n9923, new_n9924, new_n9925, new_n9926, new_n9927, new_n9928,
    new_n9929, new_n9930, new_n9931, new_n9932, new_n9933, new_n9934,
    new_n9935, new_n9936, new_n9937, new_n9938, new_n9939, new_n9940,
    new_n9941, new_n9942, new_n9943, new_n9944, new_n9945, new_n9946,
    new_n9947, new_n9948, new_n9949, new_n9950, new_n9951, new_n9952,
    new_n9953, new_n9954, new_n9955, new_n9956, new_n9957, new_n9958,
    new_n9959, new_n9960, new_n9961, new_n9962, new_n9963, new_n9964,
    new_n9965, new_n9966, new_n9967, new_n9968, new_n9969, new_n9970,
    new_n9971, new_n9972, new_n9973, new_n9974, new_n9975, new_n9976,
    new_n9977, new_n9978, new_n9979, new_n9980, new_n9981, new_n9982,
    new_n9983, new_n9984, new_n9985, new_n9986, new_n9987, new_n9988,
    new_n9989, new_n9990, new_n9991, new_n9992, new_n9993, new_n9994,
    new_n9995, new_n9996, new_n9997, new_n9998, new_n9999, new_n10000,
    new_n10001, new_n10002, new_n10003, new_n10004, new_n10005, new_n10006,
    new_n10007, new_n10008, new_n10009, new_n10010, new_n10011, new_n10012,
    new_n10013, new_n10014, new_n10015, new_n10016, new_n10017, new_n10018,
    new_n10019, new_n10020, new_n10021, new_n10022, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173, new_n10174,
    new_n10175, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180,
    new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186,
    new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192,
    new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198,
    new_n10199, new_n10200, new_n10201, new_n10202, new_n10203, new_n10204,
    new_n10205, new_n10206, new_n10207, new_n10208, new_n10209, new_n10210,
    new_n10211, new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217, new_n10218, new_n10219, new_n10220, new_n10221, new_n10222,
    new_n10223, new_n10224, new_n10225, new_n10226, new_n10227, new_n10228,
    new_n10229, new_n10230, new_n10231, new_n10232, new_n10233, new_n10234,
    new_n10235, new_n10236, new_n10237, new_n10238, new_n10239, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244, new_n10245, new_n10246,
    new_n10247, new_n10248, new_n10249, new_n10250, new_n10251, new_n10252,
    new_n10253, new_n10254, new_n10255, new_n10256, new_n10257, new_n10258,
    new_n10259, new_n10260, new_n10261, new_n10262, new_n10263, new_n10264,
    new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270,
    new_n10271, new_n10272, new_n10273, new_n10274, new_n10275, new_n10276,
    new_n10277, new_n10278, new_n10279, new_n10280, new_n10281, new_n10282,
    new_n10283, new_n10284, new_n10285, new_n10286, new_n10287, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300,
    new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306,
    new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312,
    new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318,
    new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326, new_n10327, new_n10328, new_n10329, new_n10330,
    new_n10331, new_n10332, new_n10333, new_n10334, new_n10335, new_n10336,
    new_n10337, new_n10338, new_n10339, new_n10340, new_n10341, new_n10342,
    new_n10343, new_n10344, new_n10345, new_n10346, new_n10347, new_n10348,
    new_n10349, new_n10350, new_n10351, new_n10352, new_n10353, new_n10354,
    new_n10355, new_n10356, new_n10357, new_n10358, new_n10359, new_n10360,
    new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366,
    new_n10367, new_n10368, new_n10369, new_n10370, new_n10371, new_n10372,
    new_n10373, new_n10374, new_n10375, new_n10376, new_n10377, new_n10378,
    new_n10379, new_n10380, new_n10381, new_n10382, new_n10383, new_n10384,
    new_n10385, new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391, new_n10392, new_n10393, new_n10394, new_n10395, new_n10396,
    new_n10397, new_n10398, new_n10399, new_n10400, new_n10401, new_n10402,
    new_n10403, new_n10404, new_n10405, new_n10406, new_n10407, new_n10408,
    new_n10409, new_n10410, new_n10411, new_n10412, new_n10413, new_n10414,
    new_n10415, new_n10416, new_n10417, new_n10418, new_n10419, new_n10420,
    new_n10421, new_n10422, new_n10423, new_n10424, new_n10425, new_n10426,
    new_n10427, new_n10428, new_n10429, new_n10430, new_n10431, new_n10432,
    new_n10433, new_n10434, new_n10435, new_n10436, new_n10437, new_n10438,
    new_n10439, new_n10440, new_n10441, new_n10442, new_n10443, new_n10444,
    new_n10445, new_n10446, new_n10447, new_n10448, new_n10449, new_n10450,
    new_n10451, new_n10452, new_n10453, new_n10454, new_n10455, new_n10456,
    new_n10457, new_n10458, new_n10459, new_n10460, new_n10461, new_n10462,
    new_n10463, new_n10464, new_n10465, new_n10466, new_n10467, new_n10468,
    new_n10469, new_n10470, new_n10471, new_n10472, new_n10473, new_n10474,
    new_n10475, new_n10476, new_n10477, new_n10478, new_n10479, new_n10480,
    new_n10481, new_n10482, new_n10483, new_n10484, new_n10485, new_n10486,
    new_n10487, new_n10488, new_n10489, new_n10490, new_n10491, new_n10492,
    new_n10493, new_n10494, new_n10495, new_n10496, new_n10497, new_n10498,
    new_n10499, new_n10500, new_n10501, new_n10502, new_n10503, new_n10504,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510,
    new_n10511, new_n10512, new_n10513, new_n10514, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525, new_n10526, new_n10527, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539, new_n10540,
    new_n10541, new_n10542, new_n10543, new_n10544, new_n10545, new_n10546,
    new_n10547, new_n10548, new_n10549, new_n10550, new_n10551, new_n10552,
    new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558,
    new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564,
    new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570,
    new_n10571, new_n10572, new_n10573, new_n10574, new_n10575, new_n10576,
    new_n10577, new_n10578, new_n10579, new_n10580, new_n10581, new_n10582,
    new_n10583, new_n10584, new_n10585, new_n10586, new_n10587, new_n10588,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593, new_n10594,
    new_n10595, new_n10596, new_n10597, new_n10598, new_n10599, new_n10600,
    new_n10601, new_n10602, new_n10603, new_n10604, new_n10605, new_n10606,
    new_n10607, new_n10608, new_n10609, new_n10610, new_n10611, new_n10612,
    new_n10613, new_n10614, new_n10615, new_n10616, new_n10617, new_n10618,
    new_n10619, new_n10620, new_n10621, new_n10622, new_n10623, new_n10624,
    new_n10625, new_n10626, new_n10627, new_n10628, new_n10629, new_n10630,
    new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636,
    new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642,
    new_n10643, new_n10644, new_n10645, new_n10646, new_n10647, new_n10648,
    new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654,
    new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10676, new_n10677, new_n10678,
    new_n10679, new_n10680, new_n10681, new_n10682, new_n10683, new_n10684,
    new_n10685, new_n10686, new_n10687, new_n10688, new_n10689, new_n10690,
    new_n10691, new_n10692, new_n10693, new_n10694, new_n10695, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924,
    new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005, new_n11006, new_n11007, new_n11008,
    new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11074,
    new_n11075, new_n11076, new_n11077, new_n11078, new_n11079, new_n11080,
    new_n11081, new_n11082, new_n11083, new_n11084, new_n11085, new_n11086,
    new_n11087, new_n11088, new_n11089, new_n11090, new_n11091, new_n11092,
    new_n11093, new_n11094, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101, new_n11102, new_n11103, new_n11104,
    new_n11105, new_n11106, new_n11107, new_n11108, new_n11109, new_n11110,
    new_n11111, new_n11112, new_n11113, new_n11114, new_n11115, new_n11116,
    new_n11117, new_n11118, new_n11119, new_n11120, new_n11121, new_n11122,
    new_n11123, new_n11124, new_n11125, new_n11126, new_n11127, new_n11128,
    new_n11129, new_n11130, new_n11131, new_n11132, new_n11133, new_n11134,
    new_n11135, new_n11136, new_n11137, new_n11138, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11146,
    new_n11147, new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153, new_n11154, new_n11155, new_n11156, new_n11157, new_n11158,
    new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164,
    new_n11165, new_n11166, new_n11167, new_n11168, new_n11169, new_n11170,
    new_n11171, new_n11172, new_n11173, new_n11174, new_n11175, new_n11176,
    new_n11177, new_n11178, new_n11179, new_n11180, new_n11181, new_n11182,
    new_n11183, new_n11184, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192, new_n11193, new_n11194,
    new_n11195, new_n11196, new_n11197, new_n11198, new_n11199, new_n11200,
    new_n11201, new_n11202, new_n11203, new_n11204, new_n11205, new_n11206,
    new_n11207, new_n11208, new_n11209, new_n11210, new_n11211, new_n11212,
    new_n11213, new_n11214, new_n11215, new_n11216, new_n11217, new_n11218,
    new_n11219, new_n11220, new_n11221, new_n11222, new_n11223, new_n11224,
    new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230,
    new_n11231, new_n11232, new_n11233, new_n11234, new_n11235, new_n11236,
    new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242,
    new_n11243, new_n11244, new_n11245, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254,
    new_n11255, new_n11256, new_n11257, new_n11258, new_n11259, new_n11260,
    new_n11261, new_n11262, new_n11263, new_n11264, new_n11265, new_n11266,
    new_n11267, new_n11268, new_n11269, new_n11270, new_n11271, new_n11272,
    new_n11273, new_n11274, new_n11275, new_n11276, new_n11277, new_n11278,
    new_n11279, new_n11280, new_n11281, new_n11282, new_n11283, new_n11284,
    new_n11285, new_n11286, new_n11287, new_n11288, new_n11289, new_n11290,
    new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311, new_n11312, new_n11313, new_n11314,
    new_n11315, new_n11316, new_n11317, new_n11318, new_n11319, new_n11320,
    new_n11321, new_n11322, new_n11323, new_n11324, new_n11325, new_n11326,
    new_n11327, new_n11328, new_n11329, new_n11330, new_n11331, new_n11332,
    new_n11333, new_n11334, new_n11335, new_n11336, new_n11337, new_n11338,
    new_n11339, new_n11340, new_n11341, new_n11342, new_n11343, new_n11344,
    new_n11345, new_n11346, new_n11347, new_n11348, new_n11349, new_n11350,
    new_n11351, new_n11352, new_n11353, new_n11354, new_n11355, new_n11356,
    new_n11357, new_n11358, new_n11359, new_n11360, new_n11361, new_n11362,
    new_n11363, new_n11364, new_n11365, new_n11366, new_n11367, new_n11368,
    new_n11369, new_n11370, new_n11371, new_n11372, new_n11373, new_n11374,
    new_n11375, new_n11376, new_n11377, new_n11378, new_n11379, new_n11380,
    new_n11381, new_n11382, new_n11383, new_n11384, new_n11385, new_n11386,
    new_n11387, new_n11388, new_n11389, new_n11390, new_n11391, new_n11392,
    new_n11393, new_n11394, new_n11395, new_n11396, new_n11397, new_n11398,
    new_n11399, new_n11400, new_n11401, new_n11402, new_n11403, new_n11404,
    new_n11405, new_n11406, new_n11407, new_n11408, new_n11409, new_n11410,
    new_n11411, new_n11412, new_n11413, new_n11414, new_n11415, new_n11416,
    new_n11417, new_n11418, new_n11419, new_n11420, new_n11421, new_n11422,
    new_n11423, new_n11424, new_n11425, new_n11426, new_n11427, new_n11428,
    new_n11429, new_n11430, new_n11431, new_n11432, new_n11433, new_n11434,
    new_n11435, new_n11436, new_n11437, new_n11438, new_n11439, new_n11440,
    new_n11441, new_n11442, new_n11443, new_n11444, new_n11445, new_n11446,
    new_n11447, new_n11448, new_n11449, new_n11450, new_n11451, new_n11452,
    new_n11453, new_n11454, new_n11455, new_n11456, new_n11457, new_n11458,
    new_n11459, new_n11460, new_n11461, new_n11462, new_n11463, new_n11464,
    new_n11465, new_n11466, new_n11467, new_n11468, new_n11469, new_n11470,
    new_n11471, new_n11472, new_n11473, new_n11474, new_n11475, new_n11476,
    new_n11477, new_n11478, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535, new_n11536,
    new_n11537, new_n11538, new_n11539, new_n11540, new_n11541, new_n11542,
    new_n11543, new_n11544, new_n11545, new_n11546, new_n11547, new_n11548,
    new_n11549, new_n11550, new_n11551, new_n11552, new_n11553, new_n11554,
    new_n11555, new_n11556, new_n11557, new_n11558, new_n11559, new_n11560,
    new_n11561, new_n11562, new_n11563, new_n11564, new_n11565, new_n11566,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584,
    new_n11585, new_n11586, new_n11587, new_n11588, new_n11589, new_n11590,
    new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596,
    new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602,
    new_n11603, new_n11604, new_n11605, new_n11606, new_n11607, new_n11608,
    new_n11609, new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615, new_n11616, new_n11617, new_n11618, new_n11619, new_n11620,
    new_n11621, new_n11622, new_n11623, new_n11624, new_n11625, new_n11626,
    new_n11627, new_n11628, new_n11629, new_n11630, new_n11631, new_n11632,
    new_n11633, new_n11634, new_n11635, new_n11636, new_n11637, new_n11638,
    new_n11639, new_n11640, new_n11641, new_n11642, new_n11643, new_n11644,
    new_n11645, new_n11646, new_n11647, new_n11648, new_n11649, new_n11650,
    new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656,
    new_n11657, new_n11658, new_n11659, new_n11660, new_n11661, new_n11662,
    new_n11663, new_n11664, new_n11665, new_n11666, new_n11667, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673, new_n11674,
    new_n11675, new_n11676, new_n11677, new_n11678, new_n11679, new_n11680,
    new_n11681, new_n11682, new_n11683, new_n11684, new_n11685, new_n11686,
    new_n11687, new_n11688, new_n11689, new_n11690, new_n11691, new_n11692,
    new_n11693, new_n11694, new_n11695, new_n11696, new_n11697, new_n11698,
    new_n11699, new_n11700, new_n11701, new_n11702, new_n11703, new_n11704,
    new_n11705, new_n11706, new_n11707, new_n11708, new_n11709, new_n11710,
    new_n11711, new_n11712, new_n11713, new_n11714, new_n11715, new_n11716,
    new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722,
    new_n11723, new_n11724, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755, new_n11756, new_n11757, new_n11758,
    new_n11759, new_n11760, new_n11761, new_n11762, new_n11763, new_n11764,
    new_n11765, new_n11766, new_n11767, new_n11768, new_n11769, new_n11770,
    new_n11771, new_n11772, new_n11773, new_n11774, new_n11775, new_n11776,
    new_n11777, new_n11778, new_n11779, new_n11780, new_n11781, new_n11782,
    new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788,
    new_n11789, new_n11790, new_n11791, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11817, new_n11818,
    new_n11819, new_n11820, new_n11821, new_n11822, new_n11823, new_n11824,
    new_n11825, new_n11826, new_n11827, new_n11828, new_n11829, new_n11830,
    new_n11831, new_n11832, new_n11833, new_n11834, new_n11835, new_n11836,
    new_n11837, new_n11838, new_n11839, new_n11840, new_n11841, new_n11842,
    new_n11843, new_n11844, new_n11845, new_n11846, new_n11847, new_n11848,
    new_n11849, new_n11850, new_n11851, new_n11852, new_n11853, new_n11854,
    new_n11855, new_n11856, new_n11857, new_n11858, new_n11859, new_n11860,
    new_n11861, new_n11862, new_n11863, new_n11864, new_n11865, new_n11866,
    new_n11867, new_n11868, new_n11869, new_n11870, new_n11871, new_n11872,
    new_n11873, new_n11874, new_n11875, new_n11876, new_n11877, new_n11878,
    new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884,
    new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891, new_n11892, new_n11893, new_n11894, new_n11895, new_n11896,
    new_n11897, new_n11898, new_n11899, new_n11900, new_n11901, new_n11902,
    new_n11903, new_n11904, new_n11905, new_n11906, new_n11907, new_n11908,
    new_n11909, new_n11910, new_n11911, new_n11912, new_n11913, new_n11914,
    new_n11915, new_n11916, new_n11917, new_n11918, new_n11919, new_n11920,
    new_n11921, new_n11922, new_n11923, new_n11924, new_n11925, new_n11926,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956,
    new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962,
    new_n11963, new_n11964, new_n11965, new_n11966, new_n11967, new_n11968,
    new_n11969, new_n11970, new_n11971, new_n11972, new_n11973, new_n11974,
    new_n11975, new_n11976, new_n11977, new_n11978, new_n11979, new_n11980,
    new_n11981, new_n11982, new_n11983, new_n11984, new_n11985, new_n11986,
    new_n11987, new_n11988, new_n11989, new_n11990, new_n11991, new_n11992,
    new_n11993, new_n11994, new_n11995, new_n11996, new_n11997, new_n11998,
    new_n11999, new_n12000, new_n12001, new_n12002, new_n12003, new_n12004,
    new_n12005, new_n12006, new_n12007, new_n12008, new_n12009, new_n12010,
    new_n12011, new_n12012, new_n12013, new_n12014, new_n12015, new_n12016,
    new_n12017, new_n12018, new_n12019, new_n12020, new_n12021, new_n12022,
    new_n12023, new_n12024, new_n12025, new_n12026, new_n12027, new_n12028,
    new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044, new_n12045, new_n12046,
    new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052,
    new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058,
    new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064,
    new_n12065, new_n12066, new_n12067, new_n12068, new_n12069, new_n12070,
    new_n12071, new_n12072, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12108, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113, new_n12114, new_n12115, new_n12116, new_n12117, new_n12118,
    new_n12119, new_n12120, new_n12121, new_n12122, new_n12123, new_n12124,
    new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131, new_n12132, new_n12133, new_n12134, new_n12135, new_n12136,
    new_n12137, new_n12138, new_n12139, new_n12140, new_n12141, new_n12142,
    new_n12143, new_n12144, new_n12145, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221, new_n12222, new_n12223, new_n12224, new_n12225, new_n12226,
    new_n12227, new_n12228, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235, new_n12236, new_n12237, new_n12238,
    new_n12239, new_n12240, new_n12241, new_n12242, new_n12243, new_n12244,
    new_n12245, new_n12246, new_n12247, new_n12248, new_n12249, new_n12250,
    new_n12251, new_n12252, new_n12253, new_n12254, new_n12255, new_n12256,
    new_n12257, new_n12258, new_n12259, new_n12260, new_n12261, new_n12262,
    new_n12263, new_n12264, new_n12265, new_n12266, new_n12267, new_n12268,
    new_n12269, new_n12270, new_n12271, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299, new_n12300, new_n12301, new_n12302, new_n12303, new_n12304,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316,
    new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341, new_n12342, new_n12343, new_n12344, new_n12345, new_n12346,
    new_n12347, new_n12348, new_n12349, new_n12350, new_n12351, new_n12352,
    new_n12353, new_n12354, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370,
    new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382,
    new_n12383, new_n12384, new_n12385, new_n12386, new_n12387, new_n12388,
    new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394,
    new_n12395, new_n12396, new_n12397, new_n12398, new_n12399, new_n12400,
    new_n12401, new_n12402, new_n12403, new_n12404, new_n12405, new_n12406,
    new_n12407, new_n12408, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490,
    new_n12491, new_n12492, new_n12493, new_n12494, new_n12495, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507, new_n12508,
    new_n12509, new_n12510, new_n12511, new_n12512, new_n12513, new_n12514,
    new_n12515, new_n12516, new_n12517, new_n12518, new_n12519, new_n12520,
    new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526,
    new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544,
    new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550,
    new_n12551, new_n12552, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561, new_n12562,
    new_n12563, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591, new_n12592,
    new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598,
    new_n12599, new_n12600, new_n12601, new_n12602, new_n12603, new_n12604,
    new_n12605, new_n12606, new_n12607, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620, new_n12621, new_n12622,
    new_n12623, new_n12624, new_n12625, new_n12626, new_n12627, new_n12628,
    new_n12629, new_n12630, new_n12631, new_n12632, new_n12633, new_n12634,
    new_n12635, new_n12636, new_n12637, new_n12638, new_n12639, new_n12640,
    new_n12641, new_n12642, new_n12643, new_n12644, new_n12645, new_n12646,
    new_n12647, new_n12648, new_n12649, new_n12650, new_n12651, new_n12652,
    new_n12653, new_n12654, new_n12655, new_n12656, new_n12657, new_n12658,
    new_n12659, new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665, new_n12666, new_n12667, new_n12668, new_n12669, new_n12670,
    new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676,
    new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682,
    new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688,
    new_n12689, new_n12690, new_n12691, new_n12692, new_n12693, new_n12694,
    new_n12695, new_n12696, new_n12697, new_n12698, new_n12699, new_n12700,
    new_n12701, new_n12702, new_n12703, new_n12704, new_n12705, new_n12706,
    new_n12707, new_n12708, new_n12709, new_n12710, new_n12711, new_n12712,
    new_n12713, new_n12714, new_n12715, new_n12716, new_n12717, new_n12718,
    new_n12719, new_n12720, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12740, new_n12741, new_n12742,
    new_n12743, new_n12744, new_n12745, new_n12746, new_n12747, new_n12748,
    new_n12749, new_n12750, new_n12751, new_n12752, new_n12753, new_n12754,
    new_n12755, new_n12756, new_n12757, new_n12758, new_n12759, new_n12760,
    new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766,
    new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772,
    new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807, new_n12808,
    new_n12809, new_n12810, new_n12811, new_n12812, new_n12813, new_n12814,
    new_n12815, new_n12816, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821, new_n12822, new_n12823, new_n12824, new_n12825, new_n12826,
    new_n12827, new_n12828, new_n12829, new_n12830, new_n12831, new_n12832,
    new_n12833, new_n12834, new_n12835, new_n12836, new_n12837, new_n12838,
    new_n12839, new_n12840, new_n12841, new_n12842, new_n12843, new_n12844,
    new_n12845, new_n12846, new_n12847, new_n12848, new_n12849, new_n12850,
    new_n12851, new_n12852, new_n12853, new_n12854, new_n12855, new_n12856,
    new_n12857, new_n12858, new_n12859, new_n12860, new_n12861, new_n12862,
    new_n12863, new_n12864, new_n12865, new_n12866, new_n12867, new_n12868,
    new_n12869, new_n12870, new_n12871, new_n12872, new_n12873, new_n12874,
    new_n12875, new_n12876, new_n12877, new_n12878, new_n12879, new_n12880,
    new_n12881, new_n12882, new_n12883, new_n12884, new_n12885, new_n12886,
    new_n12887, new_n12888, new_n12889, new_n12890, new_n12891, new_n12892,
    new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898,
    new_n12899, new_n12900, new_n12901, new_n12902, new_n12903, new_n12904,
    new_n12905, new_n12906, new_n12907, new_n12908, new_n12909, new_n12910,
    new_n12911, new_n12912, new_n12913, new_n12914, new_n12915, new_n12916,
    new_n12917, new_n12918, new_n12919, new_n12920, new_n12921, new_n12922,
    new_n12923, new_n12924, new_n12925, new_n12926, new_n12927, new_n12928,
    new_n12929, new_n12930, new_n12931, new_n12932, new_n12933, new_n12934,
    new_n12935, new_n12936, new_n12937, new_n12938, new_n12939, new_n12940,
    new_n12941, new_n12942, new_n12943, new_n12944, new_n12945, new_n12946,
    new_n12947, new_n12948, new_n12949, new_n12950, new_n12951, new_n12952,
    new_n12953, new_n12954, new_n12955, new_n12956, new_n12957, new_n12958,
    new_n12959, new_n12960, new_n12961, new_n12962, new_n12963, new_n12964,
    new_n12965, new_n12966, new_n12967, new_n12968, new_n12969, new_n12970,
    new_n12971, new_n12972, new_n12973, new_n12974, new_n12975, new_n12976,
    new_n12977, new_n12978, new_n12979, new_n12980, new_n12981, new_n12982,
    new_n12983, new_n12984, new_n12985, new_n12986, new_n12987, new_n12988,
    new_n12989, new_n12990, new_n12991, new_n12992, new_n12993, new_n12994,
    new_n12995, new_n12996, new_n12997, new_n12998, new_n12999, new_n13000,
    new_n13001, new_n13002, new_n13003, new_n13004, new_n13005, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026, new_n13027, new_n13028, new_n13029, new_n13030,
    new_n13031, new_n13032, new_n13033, new_n13034, new_n13035, new_n13036,
    new_n13037, new_n13038, new_n13039, new_n13040, new_n13041, new_n13042,
    new_n13043, new_n13044, new_n13045, new_n13046, new_n13047, new_n13048,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053, new_n13054,
    new_n13055, new_n13056, new_n13057, new_n13058, new_n13059, new_n13060,
    new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066,
    new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072,
    new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084,
    new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090,
    new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122, new_n13123, new_n13124, new_n13125, new_n13126,
    new_n13127, new_n13128, new_n13129, new_n13130, new_n13131, new_n13132,
    new_n13133, new_n13134, new_n13135, new_n13136, new_n13137, new_n13138,
    new_n13139, new_n13140, new_n13141, new_n13142, new_n13143, new_n13144,
    new_n13145, new_n13146, new_n13147, new_n13148, new_n13149, new_n13150,
    new_n13151, new_n13152, new_n13153, new_n13154, new_n13155, new_n13156,
    new_n13157, new_n13158, new_n13159, new_n13160, new_n13161, new_n13162,
    new_n13163, new_n13164, new_n13165, new_n13166, new_n13167, new_n13168,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186,
    new_n13187, new_n13188, new_n13189, new_n13190, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198,
    new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210,
    new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13216,
    new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222,
    new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228,
    new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234,
    new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240,
    new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252,
    new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258,
    new_n13259, new_n13260, new_n13261, new_n13262, new_n13263, new_n13264,
    new_n13265, new_n13266, new_n13267, new_n13268, new_n13269, new_n13270,
    new_n13271, new_n13272, new_n13273, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294,
    new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312,
    new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318,
    new_n13319, new_n13320, new_n13321, new_n13322, new_n13323, new_n13324,
    new_n13325, new_n13326, new_n13327, new_n13328, new_n13329, new_n13330,
    new_n13331, new_n13332, new_n13333, new_n13334, new_n13335, new_n13336,
    new_n13337, new_n13338, new_n13339, new_n13340, new_n13341, new_n13342,
    new_n13343, new_n13344, new_n13345, new_n13346, new_n13347, new_n13348,
    new_n13349, new_n13350, new_n13351, new_n13352, new_n13353, new_n13354,
    new_n13355, new_n13356, new_n13357, new_n13358, new_n13359, new_n13360,
    new_n13361, new_n13362, new_n13363, new_n13364, new_n13365, new_n13366,
    new_n13367, new_n13368, new_n13369, new_n13370, new_n13371, new_n13372,
    new_n13373, new_n13374, new_n13375, new_n13376, new_n13377, new_n13378,
    new_n13379, new_n13380, new_n13381, new_n13382, new_n13383, new_n13384,
    new_n13385, new_n13386, new_n13387, new_n13388, new_n13389, new_n13390,
    new_n13391, new_n13392, new_n13393, new_n13394, new_n13395, new_n13396,
    new_n13397, new_n13398, new_n13399, new_n13400, new_n13401, new_n13402,
    new_n13403, new_n13404, new_n13405, new_n13406, new_n13407, new_n13408,
    new_n13409, new_n13410, new_n13411, new_n13412, new_n13413, new_n13414,
    new_n13415, new_n13416, new_n13417, new_n13418, new_n13419, new_n13420,
    new_n13421, new_n13422, new_n13423, new_n13424, new_n13425, new_n13426,
    new_n13427, new_n13428, new_n13429, new_n13430, new_n13431, new_n13432,
    new_n13433, new_n13434, new_n13435, new_n13436, new_n13437, new_n13438,
    new_n13439, new_n13440, new_n13441, new_n13442, new_n13443, new_n13444,
    new_n13445, new_n13446, new_n13447, new_n13448, new_n13449, new_n13450,
    new_n13451, new_n13452, new_n13453, new_n13454, new_n13455, new_n13456,
    new_n13457, new_n13458, new_n13459, new_n13460, new_n13461, new_n13462,
    new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468,
    new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474,
    new_n13475, new_n13476, new_n13477, new_n13478, new_n13479, new_n13480,
    new_n13481, new_n13482, new_n13483, new_n13484, new_n13485, new_n13486,
    new_n13487, new_n13488, new_n13489, new_n13490, new_n13491, new_n13492,
    new_n13493, new_n13494, new_n13495, new_n13496, new_n13497, new_n13498,
    new_n13499, new_n13500, new_n13501, new_n13502, new_n13503, new_n13504,
    new_n13505, new_n13506, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534,
    new_n13535, new_n13536, new_n13537, new_n13538, new_n13539, new_n13540,
    new_n13541, new_n13542, new_n13543, new_n13544, new_n13545, new_n13546,
    new_n13547, new_n13548, new_n13549, new_n13550, new_n13551, new_n13552,
    new_n13553, new_n13554, new_n13555, new_n13556, new_n13557, new_n13558,
    new_n13559, new_n13560, new_n13561, new_n13562, new_n13563, new_n13564,
    new_n13565, new_n13566, new_n13567, new_n13568, new_n13569, new_n13570,
    new_n13571, new_n13572, new_n13573, new_n13574, new_n13575, new_n13576,
    new_n13577, new_n13578, new_n13579, new_n13580, new_n13581, new_n13582,
    new_n13583, new_n13584, new_n13585, new_n13586, new_n13587, new_n13588,
    new_n13589, new_n13590, new_n13591, new_n13592, new_n13593, new_n13594,
    new_n13595, new_n13596, new_n13597, new_n13598, new_n13599, new_n13600,
    new_n13601, new_n13602, new_n13603, new_n13604, new_n13605, new_n13606,
    new_n13607, new_n13608, new_n13609, new_n13610, new_n13611, new_n13612,
    new_n13613, new_n13614, new_n13615, new_n13616, new_n13617, new_n13618,
    new_n13619, new_n13620, new_n13621, new_n13622, new_n13623, new_n13624,
    new_n13625, new_n13626, new_n13627, new_n13628, new_n13629, new_n13630,
    new_n13631, new_n13632, new_n13633, new_n13634, new_n13635, new_n13636,
    new_n13637, new_n13638, new_n13639, new_n13640, new_n13641, new_n13642,
    new_n13643, new_n13644, new_n13645, new_n13646, new_n13647, new_n13648,
    new_n13649, new_n13650, new_n13651, new_n13652, new_n13653, new_n13654,
    new_n13655, new_n13656, new_n13657, new_n13658, new_n13659, new_n13660,
    new_n13661, new_n13662, new_n13663, new_n13664, new_n13665, new_n13666,
    new_n13667, new_n13668, new_n13669, new_n13670, new_n13671, new_n13672,
    new_n13673, new_n13674, new_n13675, new_n13676, new_n13677, new_n13678,
    new_n13679, new_n13680, new_n13681, new_n13682, new_n13683, new_n13684,
    new_n13685, new_n13686, new_n13687, new_n13688, new_n13689, new_n13690,
    new_n13691, new_n13692, new_n13693, new_n13694, new_n13695, new_n13696,
    new_n13697, new_n13698, new_n13699, new_n13700, new_n13701, new_n13702,
    new_n13703, new_n13704, new_n13705, new_n13706, new_n13707, new_n13708,
    new_n13709, new_n13710, new_n13711, new_n13712, new_n13713, new_n13714,
    new_n13715, new_n13716, new_n13717, new_n13718, new_n13719, new_n13720,
    new_n13721, new_n13722, new_n13723, new_n13724, new_n13725, new_n13726,
    new_n13727, new_n13728, new_n13729, new_n13730, new_n13731, new_n13732,
    new_n13733, new_n13734, new_n13735, new_n13736, new_n13737, new_n13738,
    new_n13739, new_n13740, new_n13741, new_n13742, new_n13743, new_n13744,
    new_n13745, new_n13746, new_n13747, new_n13748, new_n13749, new_n13750,
    new_n13751, new_n13752, new_n13753, new_n13754, new_n13755, new_n13756,
    new_n13757, new_n13758, new_n13759, new_n13760, new_n13761, new_n13762,
    new_n13763, new_n13764, new_n13765, new_n13766, new_n13767, new_n13768,
    new_n13769, new_n13770, new_n13771, new_n13772, new_n13773, new_n13774,
    new_n13775, new_n13776, new_n13777, new_n13778, new_n13779, new_n13780,
    new_n13781, new_n13782, new_n13783, new_n13784, new_n13785, new_n13786,
    new_n13787, new_n13788, new_n13789, new_n13790, new_n13791, new_n13792,
    new_n13793, new_n13794, new_n13795, new_n13796, new_n13797, new_n13798,
    new_n13799, new_n13800, new_n13801, new_n13802, new_n13803, new_n13804,
    new_n13805, new_n13806, new_n13807, new_n13808, new_n13809, new_n13810,
    new_n13811, new_n13812, new_n13813, new_n13814, new_n13815, new_n13816,
    new_n13817, new_n13818, new_n13819, new_n13820, new_n13821, new_n13822,
    new_n13823, new_n13824, new_n13825, new_n13826, new_n13827, new_n13828,
    new_n13829, new_n13830, new_n13831, new_n13832, new_n13833, new_n13834,
    new_n13835, new_n13836, new_n13837, new_n13838, new_n13839, new_n13840,
    new_n13841, new_n13842, new_n13843, new_n13844, new_n13845, new_n13846,
    new_n13847, new_n13848, new_n13849, new_n13850, new_n13851, new_n13852,
    new_n13853, new_n13854, new_n13855, new_n13856, new_n13857, new_n13858,
    new_n13859, new_n13860, new_n13861, new_n13862, new_n13863, new_n13864,
    new_n13865, new_n13866, new_n13867, new_n13868, new_n13869, new_n13870,
    new_n13871, new_n13872, new_n13873, new_n13874, new_n13875, new_n13876,
    new_n13877, new_n13878, new_n13879, new_n13880, new_n13881, new_n13882,
    new_n13883, new_n13884, new_n13885, new_n13886, new_n13887, new_n13888,
    new_n13889, new_n13890, new_n13891, new_n13892, new_n13893, new_n13894,
    new_n13895, new_n13896, new_n13897, new_n13898, new_n13899, new_n13900,
    new_n13901, new_n13902, new_n13903, new_n13904, new_n13905, new_n13906,
    new_n13907, new_n13908, new_n13909, new_n13910, new_n13911, new_n13912,
    new_n13913, new_n13914, new_n13915, new_n13916, new_n13917, new_n13918,
    new_n13919, new_n13920, new_n13921, new_n13922, new_n13923, new_n13924,
    new_n13925, new_n13926, new_n13927, new_n13928, new_n13929, new_n13930,
    new_n13931, new_n13932, new_n13933, new_n13934, new_n13935, new_n13936,
    new_n13937, new_n13938, new_n13939, new_n13940, new_n13941, new_n13942,
    new_n13943, new_n13944, new_n13945, new_n13946, new_n13947, new_n13948,
    new_n13949, new_n13950, new_n13951, new_n13952, new_n13953, new_n13954,
    new_n13955, new_n13956, new_n13957, new_n13958, new_n13959, new_n13960,
    new_n13961, new_n13962, new_n13963, new_n13964, new_n13965, new_n13966,
    new_n13967, new_n13968, new_n13969, new_n13970, new_n13971, new_n13972,
    new_n13973, new_n13974, new_n13975, new_n13976, new_n13977, new_n13978,
    new_n13979, new_n13980, new_n13981, new_n13982, new_n13983, new_n13984,
    new_n13985, new_n13986, new_n13987, new_n13988, new_n13989, new_n13990,
    new_n13991, new_n13992, new_n13993, new_n13994, new_n13995, new_n13996,
    new_n13997, new_n13998, new_n13999, new_n14000, new_n14001, new_n14002,
    new_n14003, new_n14004, new_n14005, new_n14006, new_n14007, new_n14008,
    new_n14009, new_n14010, new_n14011, new_n14012, new_n14013, new_n14014,
    new_n14015, new_n14016, new_n14017, new_n14018, new_n14019, new_n14020,
    new_n14021, new_n14022, new_n14023, new_n14024, new_n14025, new_n14026,
    new_n14027, new_n14028, new_n14029, new_n14030, new_n14031, new_n14032,
    new_n14033, new_n14034, new_n14035, new_n14036, new_n14037, new_n14038,
    new_n14039, new_n14040, new_n14041, new_n14042, new_n14043, new_n14044,
    new_n14045, new_n14046, new_n14047, new_n14048, new_n14049, new_n14050,
    new_n14051, new_n14052, new_n14053, new_n14054, new_n14055, new_n14056,
    new_n14057, new_n14058, new_n14059, new_n14060, new_n14061, new_n14062,
    new_n14063, new_n14064, new_n14065, new_n14066, new_n14067, new_n14068,
    new_n14069, new_n14070, new_n14071, new_n14072, new_n14073, new_n14074,
    new_n14075, new_n14076, new_n14077, new_n14078, new_n14079, new_n14080,
    new_n14081, new_n14082, new_n14083, new_n14084, new_n14085, new_n14086,
    new_n14087, new_n14088, new_n14089, new_n14090, new_n14091, new_n14092,
    new_n14093, new_n14094, new_n14095, new_n14096, new_n14097, new_n14098,
    new_n14099, new_n14100, new_n14101, new_n14102, new_n14103, new_n14104,
    new_n14105, new_n14106, new_n14107, new_n14108, new_n14109, new_n14110,
    new_n14111, new_n14112, new_n14113, new_n14114, new_n14115, new_n14116,
    new_n14117, new_n14118, new_n14119, new_n14120, new_n14121, new_n14122,
    new_n14123, new_n14124, new_n14125, new_n14126, new_n14127, new_n14128,
    new_n14129, new_n14130, new_n14131, new_n14132, new_n14133, new_n14134,
    new_n14135, new_n14136, new_n14137, new_n14138, new_n14139, new_n14140,
    new_n14141, new_n14142, new_n14143, new_n14144, new_n14145, new_n14146,
    new_n14147, new_n14148, new_n14149, new_n14150, new_n14151, new_n14152,
    new_n14153, new_n14154, new_n14155, new_n14156, new_n14157, new_n14158,
    new_n14159, new_n14160, new_n14161, new_n14162, new_n14163, new_n14164,
    new_n14165, new_n14166, new_n14167, new_n14168, new_n14169, new_n14170,
    new_n14171, new_n14172, new_n14173, new_n14174, new_n14175, new_n14176,
    new_n14177, new_n14178, new_n14179, new_n14180, new_n14181, new_n14182,
    new_n14183, new_n14184, new_n14185, new_n14186, new_n14187, new_n14188,
    new_n14189, new_n14190, new_n14191, new_n14192, new_n14193, new_n14194,
    new_n14195, new_n14196, new_n14197, new_n14198, new_n14199, new_n14200,
    new_n14201, new_n14202, new_n14203, new_n14204, new_n14205, new_n14206,
    new_n14207, new_n14208, new_n14209, new_n14210, new_n14211, new_n14212,
    new_n14213, new_n14214, new_n14215, new_n14216, new_n14217, new_n14218,
    new_n14219, new_n14220, new_n14221, new_n14222, new_n14223, new_n14224,
    new_n14225, new_n14226, new_n14227, new_n14228, new_n14229, new_n14230,
    new_n14231, new_n14232, new_n14233, new_n14234, new_n14235, new_n14236,
    new_n14237, new_n14238, new_n14239, new_n14240, new_n14241, new_n14242,
    new_n14243, new_n14244, new_n14245, new_n14246, new_n14247, new_n14248,
    new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254,
    new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260,
    new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267, new_n14268, new_n14269, new_n14270, new_n14271, new_n14272,
    new_n14273, new_n14274, new_n14275, new_n14276, new_n14277, new_n14278,
    new_n14279, new_n14280, new_n14281, new_n14282, new_n14283, new_n14284,
    new_n14285, new_n14286, new_n14287, new_n14288, new_n14289, new_n14290,
    new_n14291, new_n14292, new_n14293, new_n14294, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310, new_n14311, new_n14312, new_n14313, new_n14314,
    new_n14315, new_n14316, new_n14317, new_n14318, new_n14319, new_n14320,
    new_n14321, new_n14322, new_n14323, new_n14324, new_n14325, new_n14326,
    new_n14327, new_n14328, new_n14329, new_n14330, new_n14331, new_n14332,
    new_n14333, new_n14334, new_n14335, new_n14336, new_n14337, new_n14338,
    new_n14339, new_n14340, new_n14341, new_n14342, new_n14343, new_n14344,
    new_n14345, new_n14346, new_n14347, new_n14348, new_n14349, new_n14350,
    new_n14351, new_n14352, new_n14353, new_n14354, new_n14355, new_n14356,
    new_n14357, new_n14358, new_n14359, new_n14360, new_n14361, new_n14362,
    new_n14363, new_n14364, new_n14365, new_n14366, new_n14367, new_n14368,
    new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374,
    new_n14375, new_n14376, new_n14377, new_n14378, new_n14379, new_n14380,
    new_n14381, new_n14382, new_n14383, new_n14384, new_n14385, new_n14386,
    new_n14387, new_n14388, new_n14389, new_n14390, new_n14391, new_n14392,
    new_n14393, new_n14394, new_n14395, new_n14396, new_n14397, new_n14398,
    new_n14399, new_n14400, new_n14401, new_n14402, new_n14403, new_n14404,
    new_n14405, new_n14406, new_n14407, new_n14408, new_n14409, new_n14410,
    new_n14411, new_n14412, new_n14413, new_n14414, new_n14415, new_n14416,
    new_n14417, new_n14418, new_n14419, new_n14420, new_n14421, new_n14422,
    new_n14423, new_n14424, new_n14425, new_n14426, new_n14427, new_n14428,
    new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439, new_n14440,
    new_n14441, new_n14442, new_n14443, new_n14444, new_n14445, new_n14446,
    new_n14447, new_n14448, new_n14449, new_n14450, new_n14451, new_n14452,
    new_n14453, new_n14454, new_n14455, new_n14456, new_n14457, new_n14458,
    new_n14459, new_n14460, new_n14461, new_n14462, new_n14463, new_n14464,
    new_n14465, new_n14466, new_n14467, new_n14468, new_n14469, new_n14470,
    new_n14471, new_n14472, new_n14473, new_n14474, new_n14475, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510, new_n14511, new_n14512,
    new_n14513, new_n14514, new_n14515, new_n14516, new_n14517, new_n14518,
    new_n14519, new_n14520, new_n14521, new_n14522, new_n14523, new_n14524,
    new_n14525, new_n14526, new_n14527, new_n14528, new_n14529, new_n14530,
    new_n14531, new_n14532, new_n14533, new_n14534, new_n14535, new_n14536,
    new_n14537, new_n14538, new_n14539, new_n14540, new_n14541, new_n14542,
    new_n14543, new_n14544, new_n14545, new_n14546, new_n14547, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570, new_n14571, new_n14572,
    new_n14573, new_n14574, new_n14575, new_n14576, new_n14577, new_n14578,
    new_n14579, new_n14580, new_n14581, new_n14582, new_n14583, new_n14584,
    new_n14585, new_n14586, new_n14587, new_n14588, new_n14589, new_n14590,
    new_n14591, new_n14592, new_n14593, new_n14594, new_n14595, new_n14596,
    new_n14597, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602,
    new_n14603, new_n14604, new_n14605, new_n14606, new_n14607, new_n14608,
    new_n14609, new_n14610, new_n14611, new_n14612, new_n14613, new_n14614,
    new_n14615, new_n14616, new_n14617, new_n14618, new_n14619, new_n14620,
    new_n14621, new_n14622, new_n14623, new_n14624, new_n14625, new_n14626,
    new_n14627, new_n14628, new_n14629, new_n14630, new_n14631, new_n14632,
    new_n14633, new_n14634, new_n14635, new_n14636, new_n14637, new_n14638,
    new_n14639, new_n14640, new_n14641, new_n14642, new_n14643, new_n14644,
    new_n14645, new_n14646, new_n14647, new_n14648, new_n14649, new_n14650,
    new_n14651, new_n14652, new_n14653, new_n14654, new_n14655, new_n14656,
    new_n14657, new_n14658, new_n14659, new_n14660, new_n14661, new_n14662,
    new_n14663, new_n14664, new_n14665, new_n14666, new_n14667, new_n14668,
    new_n14669, new_n14670, new_n14671, new_n14672, new_n14673, new_n14674,
    new_n14675, new_n14676, new_n14677, new_n14678, new_n14679, new_n14680,
    new_n14681, new_n14682, new_n14683, new_n14684, new_n14685, new_n14686,
    new_n14687, new_n14688, new_n14689, new_n14690, new_n14691, new_n14692,
    new_n14693, new_n14694, new_n14695, new_n14696, new_n14697, new_n14698,
    new_n14699, new_n14700, new_n14701, new_n14702, new_n14703, new_n14704,
    new_n14705, new_n14706, new_n14707, new_n14708, new_n14709, new_n14710,
    new_n14711, new_n14712, new_n14713, new_n14714, new_n14715, new_n14716,
    new_n14717, new_n14718, new_n14719, new_n14720, new_n14721, new_n14722,
    new_n14723, new_n14724, new_n14725, new_n14726, new_n14727, new_n14728,
    new_n14729, new_n14730, new_n14731, new_n14732, new_n14733, new_n14734,
    new_n14735, new_n14736, new_n14737, new_n14738, new_n14739, new_n14740,
    new_n14741, new_n14742, new_n14743, new_n14744, new_n14745, new_n14746,
    new_n14747, new_n14748, new_n14749, new_n14750, new_n14751, new_n14752,
    new_n14753, new_n14754, new_n14755, new_n14756, new_n14757, new_n14758,
    new_n14759, new_n14760, new_n14761, new_n14762, new_n14763, new_n14764,
    new_n14765, new_n14766, new_n14767, new_n14768, new_n14769, new_n14770,
    new_n14771, new_n14772, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800,
    new_n14801, new_n14802, new_n14803, new_n14804, new_n14805, new_n14806,
    new_n14807, new_n14808, new_n14809, new_n14810, new_n14811, new_n14812,
    new_n14813, new_n14814, new_n14815, new_n14816, new_n14817, new_n14818,
    new_n14819, new_n14820, new_n14821, new_n14822, new_n14823, new_n14824,
    new_n14825, new_n14826, new_n14827, new_n14828, new_n14829, new_n14830,
    new_n14831, new_n14832, new_n14833, new_n14834, new_n14835, new_n14836,
    new_n14837, new_n14838, new_n14839, new_n14840, new_n14841, new_n14842,
    new_n14843, new_n14844, new_n14845, new_n14846, new_n14847, new_n14848,
    new_n14849, new_n14850, new_n14851, new_n14852, new_n14853, new_n14854,
    new_n14855, new_n14856, new_n14857, new_n14858, new_n14859, new_n14860,
    new_n14861, new_n14862, new_n14863, new_n14864, new_n14865, new_n14866,
    new_n14867, new_n14868, new_n14869, new_n14870, new_n14871, new_n14872,
    new_n14873, new_n14874, new_n14875, new_n14876, new_n14877, new_n14878,
    new_n14879, new_n14880, new_n14881, new_n14882, new_n14883, new_n14884,
    new_n14885, new_n14886, new_n14887, new_n14888, new_n14889, new_n14890,
    new_n14891, new_n14892, new_n14893, new_n14894, new_n14895, new_n14896,
    new_n14897, new_n14898, new_n14899, new_n14900, new_n14901, new_n14902,
    new_n14903, new_n14904, new_n14905, new_n14906, new_n14907, new_n14908,
    new_n14909, new_n14910, new_n14911, new_n14912, new_n14913, new_n14914,
    new_n14915, new_n14916, new_n14917, new_n14918, new_n14919, new_n14920,
    new_n14921, new_n14922, new_n14923, new_n14924, new_n14925, new_n14926,
    new_n14927, new_n14928, new_n14929, new_n14930, new_n14931, new_n14932,
    new_n14933, new_n14934, new_n14935, new_n14936, new_n14937, new_n14938,
    new_n14939, new_n14940, new_n14941, new_n14942, new_n14943, new_n14944,
    new_n14945, new_n14946, new_n14947, new_n14948, new_n14949, new_n14950,
    new_n14951, new_n14952, new_n14953, new_n14954, new_n14955, new_n14956,
    new_n14957, new_n14958, new_n14959, new_n14960, new_n14961, new_n14962,
    new_n14963, new_n14964, new_n14965, new_n14966, new_n14967, new_n14968,
    new_n14969, new_n14970, new_n14971, new_n14972, new_n14973, new_n14974,
    new_n14975, new_n14976, new_n14977, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986,
    new_n14987, new_n14988, new_n14989, new_n14990, new_n14991, new_n14992,
    new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998,
    new_n14999, new_n15000, new_n15001, new_n15002, new_n15003, new_n15004,
    new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011, new_n15012, new_n15013, new_n15014, new_n15015, new_n15016,
    new_n15017, new_n15018, new_n15019, new_n15020, new_n15021, new_n15022,
    new_n15023, new_n15024, new_n15025, new_n15026, new_n15027, new_n15028,
    new_n15029, new_n15030, new_n15031, new_n15032, new_n15033, new_n15034,
    new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040,
    new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046,
    new_n15047, new_n15048, new_n15049, new_n15050, new_n15051, new_n15052,
    new_n15053, new_n15054, new_n15055, new_n15056, new_n15057, new_n15058,
    new_n15059, new_n15060, new_n15061, new_n15062, new_n15063, new_n15064,
    new_n15065, new_n15066, new_n15067, new_n15068, new_n15069, new_n15070,
    new_n15071, new_n15072, new_n15073, new_n15074, new_n15075, new_n15076,
    new_n15077, new_n15078, new_n15079, new_n15080, new_n15081, new_n15082,
    new_n15083, new_n15084, new_n15085, new_n15086, new_n15087, new_n15088,
    new_n15089, new_n15090, new_n15091, new_n15092, new_n15093, new_n15094,
    new_n15095, new_n15096, new_n15097, new_n15098, new_n15099, new_n15100,
    new_n15101, new_n15102, new_n15103, new_n15104, new_n15105, new_n15106,
    new_n15107, new_n15108, new_n15109, new_n15110, new_n15111, new_n15112,
    new_n15113, new_n15114, new_n15115, new_n15116, new_n15117, new_n15118,
    new_n15119, new_n15120, new_n15121, new_n15122, new_n15123, new_n15124,
    new_n15125, new_n15126, new_n15127, new_n15128, new_n15129, new_n15130,
    new_n15131, new_n15132, new_n15133, new_n15134, new_n15135, new_n15136,
    new_n15137, new_n15138, new_n15139, new_n15140, new_n15141, new_n15142,
    new_n15143, new_n15144, new_n15145, new_n15146, new_n15147, new_n15148,
    new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154,
    new_n15155, new_n15156, new_n15157, new_n15158, new_n15159, new_n15160,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165, new_n15166,
    new_n15167, new_n15168, new_n15169, new_n15170, new_n15171, new_n15172,
    new_n15173, new_n15174, new_n15175, new_n15176, new_n15177, new_n15178,
    new_n15179, new_n15180, new_n15181, new_n15182, new_n15183, new_n15184,
    new_n15185, new_n15186, new_n15187, new_n15188, new_n15189, new_n15190,
    new_n15191, new_n15192, new_n15193, new_n15194, new_n15195, new_n15196,
    new_n15197, new_n15198, new_n15199, new_n15200, new_n15201, new_n15202,
    new_n15203, new_n15204, new_n15205, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230, new_n15231, new_n15232,
    new_n15233, new_n15234, new_n15235, new_n15236, new_n15237, new_n15238,
    new_n15239, new_n15240, new_n15241, new_n15242, new_n15243, new_n15244,
    new_n15245, new_n15246, new_n15247, new_n15248, new_n15249, new_n15250,
    new_n15251, new_n15252, new_n15253, new_n15254, new_n15255, new_n15256,
    new_n15257, new_n15258, new_n15259, new_n15260, new_n15261, new_n15262,
    new_n15263, new_n15264, new_n15265, new_n15266, new_n15267, new_n15268,
    new_n15269, new_n15270, new_n15271, new_n15272, new_n15273, new_n15274,
    new_n15275, new_n15276, new_n15277, new_n15278, new_n15279, new_n15280,
    new_n15281, new_n15282, new_n15283, new_n15284, new_n15285, new_n15286,
    new_n15287, new_n15288, new_n15289, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300, new_n15301, new_n15302, new_n15303, new_n15304,
    new_n15305, new_n15306, new_n15307, new_n15308, new_n15309, new_n15310,
    new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316,
    new_n15317, new_n15318, new_n15319, new_n15320, new_n15321, new_n15322,
    new_n15323, new_n15324, new_n15325, new_n15326, new_n15327, new_n15328,
    new_n15329, new_n15330, new_n15331, new_n15332, new_n15333, new_n15334,
    new_n15335, new_n15336, new_n15337, new_n15338, new_n15339, new_n15340,
    new_n15341, new_n15342, new_n15343, new_n15344, new_n15345, new_n15346,
    new_n15347, new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353, new_n15354, new_n15355, new_n15356, new_n15357, new_n15358,
    new_n15359, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15366, new_n15367, new_n15368, new_n15369, new_n15370,
    new_n15371, new_n15372, new_n15373, new_n15374, new_n15375, new_n15376,
    new_n15377, new_n15378, new_n15379, new_n15380, new_n15381, new_n15382,
    new_n15383, new_n15384, new_n15385, new_n15386, new_n15387, new_n15388,
    new_n15389, new_n15390, new_n15391, new_n15392, new_n15393, new_n15394,
    new_n15395, new_n15396, new_n15397, new_n15398, new_n15399, new_n15400,
    new_n15401, new_n15402, new_n15403, new_n15404, new_n15405, new_n15406,
    new_n15407, new_n15408, new_n15409, new_n15410, new_n15411, new_n15412,
    new_n15413, new_n15414, new_n15415, new_n15416, new_n15417, new_n15418,
    new_n15419, new_n15420, new_n15421, new_n15422, new_n15423, new_n15424,
    new_n15425, new_n15426, new_n15427, new_n15428, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435, new_n15436,
    new_n15437, new_n15438, new_n15439, new_n15440, new_n15441, new_n15442,
    new_n15443, new_n15444, new_n15445, new_n15446, new_n15447, new_n15448,
    new_n15449, new_n15450, new_n15451, new_n15452, new_n15453, new_n15454,
    new_n15455, new_n15456, new_n15457, new_n15458, new_n15459, new_n15460,
    new_n15461, new_n15462, new_n15463, new_n15464, new_n15465, new_n15466,
    new_n15467, new_n15468, new_n15469, new_n15470, new_n15471, new_n15472,
    new_n15473, new_n15474, new_n15475, new_n15476, new_n15477, new_n15478,
    new_n15479, new_n15480, new_n15481, new_n15482, new_n15483, new_n15484,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489, new_n15490,
    new_n15491, new_n15492, new_n15493, new_n15494, new_n15495, new_n15496,
    new_n15497, new_n15498, new_n15499, new_n15500, new_n15501, new_n15502,
    new_n15503, new_n15504, new_n15505, new_n15506, new_n15507, new_n15508,
    new_n15509, new_n15510, new_n15511, new_n15512, new_n15513, new_n15514,
    new_n15515, new_n15516, new_n15517, new_n15518, new_n15519, new_n15520,
    new_n15521, new_n15522, new_n15523, new_n15524, new_n15525, new_n15526,
    new_n15527, new_n15528, new_n15529, new_n15530, new_n15531, new_n15532,
    new_n15533, new_n15534, new_n15535, new_n15536, new_n15537, new_n15538,
    new_n15539, new_n15540, new_n15541, new_n15542, new_n15543, new_n15544,
    new_n15545, new_n15546, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555, new_n15556,
    new_n15557, new_n15558, new_n15559, new_n15560, new_n15561, new_n15562,
    new_n15563, new_n15564, new_n15565, new_n15566, new_n15567, new_n15568,
    new_n15569, new_n15570, new_n15571, new_n15572, new_n15573, new_n15574,
    new_n15575, new_n15576, new_n15577, new_n15578, new_n15579, new_n15580,
    new_n15581, new_n15582, new_n15583, new_n15584, new_n15585, new_n15586,
    new_n15587, new_n15588, new_n15589, new_n15590, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597, new_n15598,
    new_n15599, new_n15600, new_n15601, new_n15602, new_n15603, new_n15604,
    new_n15605, new_n15606, new_n15607, new_n15608, new_n15609, new_n15610,
    new_n15611, new_n15612, new_n15613, new_n15614, new_n15615, new_n15616,
    new_n15617, new_n15618, new_n15619, new_n15620, new_n15621, new_n15622,
    new_n15623, new_n15624, new_n15625, new_n15626, new_n15627, new_n15628,
    new_n15629, new_n15630, new_n15631, new_n15632, new_n15633, new_n15634,
    new_n15635, new_n15636, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646,
    new_n15647, new_n15648, new_n15649, new_n15650, new_n15651, new_n15652,
    new_n15653, new_n15654, new_n15655, new_n15656, new_n15657, new_n15658,
    new_n15659, new_n15660, new_n15661, new_n15662, new_n15663, new_n15664,
    new_n15665, new_n15666, new_n15667, new_n15668, new_n15669, new_n15670,
    new_n15671, new_n15672, new_n15673, new_n15674, new_n15675, new_n15676,
    new_n15677, new_n15678, new_n15679, new_n15680, new_n15681, new_n15682,
    new_n15683, new_n15684, new_n15685, new_n15686, new_n15687, new_n15688,
    new_n15689, new_n15690, new_n15691, new_n15692, new_n15693, new_n15694,
    new_n15695, new_n15696, new_n15697, new_n15698, new_n15699, new_n15700,
    new_n15701, new_n15702, new_n15703, new_n15704, new_n15705, new_n15706,
    new_n15707, new_n15708, new_n15709, new_n15710, new_n15711, new_n15712,
    new_n15713, new_n15714, new_n15715, new_n15716, new_n15717, new_n15718,
    new_n15719, new_n15720, new_n15721, new_n15722, new_n15723, new_n15724,
    new_n15725, new_n15726, new_n15727, new_n15728, new_n15729, new_n15730,
    new_n15731, new_n15732, new_n15733, new_n15734, new_n15735, new_n15736,
    new_n15737, new_n15738, new_n15739, new_n15740, new_n15741, new_n15742,
    new_n15743, new_n15744, new_n15745, new_n15746, new_n15747, new_n15748,
    new_n15749, new_n15750, new_n15751, new_n15752, new_n15753, new_n15754,
    new_n15755, new_n15756, new_n15757, new_n15758, new_n15759, new_n15760,
    new_n15761, new_n15762, new_n15763, new_n15764, new_n15765, new_n15766,
    new_n15767, new_n15768, new_n15769, new_n15770, new_n15771, new_n15772,
    new_n15773, new_n15774, new_n15775, new_n15776, new_n15777, new_n15778,
    new_n15779, new_n15780, new_n15781, new_n15782, new_n15783, new_n15784,
    new_n15785, new_n15786, new_n15787, new_n15788, new_n15789, new_n15790,
    new_n15791, new_n15792, new_n15793, new_n15794, new_n15795, new_n15796,
    new_n15797, new_n15798, new_n15799, new_n15800, new_n15801, new_n15802,
    new_n15803, new_n15804, new_n15805, new_n15806, new_n15807, new_n15808,
    new_n15809, new_n15810, new_n15811, new_n15812, new_n15813, new_n15814,
    new_n15815, new_n15816, new_n15817, new_n15818, new_n15819, new_n15820,
    new_n15821, new_n15822, new_n15823, new_n15824, new_n15825, new_n15826,
    new_n15827, new_n15828, new_n15829, new_n15830, new_n15831, new_n15832,
    new_n15833, new_n15834, new_n15835, new_n15836, new_n15837, new_n15838,
    new_n15839, new_n15840, new_n15841, new_n15842, new_n15843, new_n15844,
    new_n15845, new_n15846, new_n15847, new_n15848, new_n15849, new_n15850,
    new_n15851, new_n15852, new_n15853, new_n15854, new_n15855, new_n15856,
    new_n15857, new_n15858, new_n15859, new_n15860, new_n15861, new_n15862,
    new_n15863, new_n15864, new_n15865, new_n15866, new_n15867, new_n15868,
    new_n15869, new_n15870, new_n15871, new_n15872, new_n15873, new_n15874,
    new_n15875, new_n15876, new_n15877, new_n15878, new_n15879, new_n15880,
    new_n15881, new_n15882, new_n15883, new_n15884, new_n15885, new_n15886,
    new_n15887, new_n15888, new_n15889, new_n15890, new_n15891, new_n15892,
    new_n15893, new_n15894, new_n15895, new_n15896, new_n15897, new_n15898,
    new_n15899, new_n15900, new_n15901, new_n15902, new_n15903, new_n15904,
    new_n15905, new_n15906, new_n15907, new_n15908, new_n15909, new_n15910,
    new_n15911, new_n15912, new_n15913, new_n15914, new_n15915, new_n15916,
    new_n15917, new_n15918, new_n15919, new_n15920, new_n15921, new_n15922,
    new_n15923, new_n15924, new_n15925, new_n15926, new_n15927, new_n15928,
    new_n15929, new_n15930, new_n15931, new_n15932, new_n15933, new_n15934,
    new_n15935, new_n15936, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947, new_n15948, new_n15949, new_n15950, new_n15951, new_n15952,
    new_n15953, new_n15954;
  assign new_n4097 = n2022 ^ n2020;
  assign new_n4098 = ~n2020 & n2021;
  assign new_n4099 = new_n4098 ^ n2020;
  assign new_n4100 = new_n4099 ^ n2021;
  assign new_n4101 = ~n2022 & new_n4100;
  assign new_n4102 = new_n4101 ^ new_n4100;
  assign new_n4103 = n2021 & n2022;
  assign new_n4104 = new_n4103 ^ n2020;
  assign new_n4105 = new_n4104 ^ new_n4102;
  assign new_n4106 = new_n4105 ^ new_n4097;
  assign new_n4107 = new_n4106 ^ new_n4099;
  assign new_n4108 = ~n2044 & ~n2045;
  assign new_n4109 = n2043 & new_n4108;
  assign new_n4110 = new_n4109 ^ new_n4108;
  assign new_n4111 = ~new_n4107 & new_n4110;
  assign new_n4112 = ~n2046 & ~n2047;
  assign new_n4113 = ~n2048 & new_n4112;
  assign new_n4114 = new_n4113 ^ new_n4112;
  assign new_n4115 = new_n4114 ^ n2046;
  assign new_n4116 = ~n2017 & ~n2019;
  assign new_n4117 = n2018 & new_n4116;
  assign new_n4118 = new_n4117 ^ new_n4116;
  assign new_n4119 = ~new_n4115 & new_n4118;
  assign new_n4120 = new_n4111 & new_n4119;
  assign new_n4121 = n2038 & new_n4120;
  assign new_n4122 = n2039 & new_n4120;
  assign new_n4123 = n2040 & new_n4120;
  assign new_n4124 = n2042 & new_n4120;
  assign new_n4125 = n2041 & new_n4120;
  assign new_n4126 = new_n4124 & new_n4125;
  assign new_n4127 = new_n4124 ^ n2041;
  assign new_n4128 = new_n4127 ^ new_n4126;
  assign new_n4129 = n2017 & n2018;
  assign new_n4130 = new_n4129 ^ n2017;
  assign new_n4131 = new_n4130 ^ n2018;
  assign new_n4132 = new_n4131 ^ new_n4118;
  assign new_n4133 = ~new_n4132 & new_n4104;
  assign new_n4134 = new_n4133 ^ new_n4132;
  assign new_n4135 = ~n2022 & new_n4098;
  assign new_n4136 = new_n4135 ^ new_n4098;
  assign new_n4137 = new_n4136 ^ new_n4103;
  assign new_n4138 = ~new_n4132 & new_n4137;
  assign new_n4139 = new_n4138 ^ new_n4134;
  assign new_n4140 = n2019 & new_n4130;
  assign new_n4141 = ~new_n4099 & new_n4140;
  assign new_n4142 = new_n4140 ^ new_n4130;
  assign new_n4143 = ~n2021 & new_n4142;
  assign new_n4144 = ~new_n4141 & ~new_n4143;
  assign new_n4145 = new_n4136 ^ n2022;
  assign new_n4146 = ~new_n4145 & new_n4142;
  assign new_n4147 = new_n4106 ^ n2020;
  assign new_n4148 = ~new_n4147 & new_n4140;
  assign new_n4149 = ~new_n4146 & ~new_n4148;
  assign new_n4150 = ~new_n4149 & new_n4144;
  assign new_n4151 = new_n4150 ^ new_n4144;
  assign new_n4152 = new_n4151 ^ new_n4139;
  assign new_n4153 = new_n4152 ^ new_n4133;
  assign new_n4154 = new_n4128 & new_n4153;
  assign new_n4155 = n2041 & new_n4153;
  assign new_n4156 = new_n4155 ^ new_n4154;
  assign new_n4157 = n2042 & new_n4153;
  assign new_n4158 = new_n4157 ^ new_n4156;
  assign new_n4159 = ~new_n4120 & new_n4157;
  assign new_n4160 = new_n4159 ^ new_n4158;
  assign new_n4161 = new_n4160 ^ new_n4124;
  assign new_n4162 = n2040 & new_n4153;
  assign new_n4163 = ~new_n4162 & new_n4124;
  assign new_n4164 = new_n4163 ^ new_n4162;
  assign new_n4165 = new_n4164 ^ new_n4161;
  assign new_n4166 = new_n4125 & new_n4164;
  assign new_n4167 = new_n4166 ^ new_n4164;
  assign new_n4168 = new_n4128 ^ n2041;
  assign new_n4169 = new_n4168 ^ new_n4125;
  assign new_n4170 = new_n4169 ^ new_n4167;
  assign new_n4171 = new_n4170 ^ new_n4165;
  assign new_n4172 = n2039 & new_n4153;
  assign new_n4173 = ~new_n4124 & ~new_n4172;
  assign new_n4174 = new_n4173 ^ new_n4172;
  assign new_n4175 = n2038 & new_n4153;
  assign new_n4176 = ~new_n4175 & new_n4124;
  assign new_n4177 = new_n4176 ^ new_n4175;
  assign new_n4178 = new_n4177 ^ new_n4174;
  assign new_n4179 = new_n4125 & new_n4178;
  assign new_n4180 = new_n4179 ^ new_n4178;
  assign new_n4181 = ~new_n4171 & ~new_n4180;
  assign new_n4182 = ~new_n4123 & ~new_n4181;
  assign new_n4183 = new_n4182 ^ new_n4181;
  assign new_n4184 = n2037 & new_n4153;
  assign new_n4185 = ~new_n4124 & ~new_n4184;
  assign new_n4186 = new_n4185 ^ new_n4184;
  assign new_n4187 = n2036 & new_n4153;
  assign new_n4188 = ~new_n4187 & new_n4124;
  assign new_n4189 = new_n4188 ^ new_n4187;
  assign new_n4190 = new_n4189 ^ new_n4186;
  assign new_n4191 = ~new_n4125 & new_n4190;
  assign new_n4192 = new_n4191 ^ new_n4190;
  assign new_n4193 = n2035 & new_n4153;
  assign new_n4194 = ~new_n4124 & ~new_n4193;
  assign new_n4195 = new_n4194 ^ new_n4193;
  assign new_n4196 = n2034 & new_n4153;
  assign new_n4197 = ~new_n4196 & new_n4124;
  assign new_n4198 = new_n4197 ^ new_n4196;
  assign new_n4199 = new_n4198 ^ new_n4195;
  assign new_n4200 = new_n4125 & new_n4199;
  assign new_n4201 = new_n4200 ^ new_n4199;
  assign new_n4202 = ~new_n4192 & ~new_n4201;
  assign new_n4203 = ~new_n4202 & new_n4123;
  assign new_n4204 = new_n4203 ^ new_n4202;
  assign new_n4205 = new_n4183 & new_n4204;
  assign new_n4206 = ~new_n4205 & new_n4122;
  assign new_n4207 = new_n4206 ^ new_n4205;
  assign new_n4208 = n2044 & new_n4153;
  assign new_n4209 = ~new_n4169 & new_n4208;
  assign new_n4210 = new_n4209 ^ new_n4124;
  assign new_n4211 = ~new_n4208 & new_n4124;
  assign new_n4212 = new_n4211 ^ new_n4208;
  assign new_n4213 = new_n4212 ^ new_n4210;
  assign new_n4214 = new_n4213 ^ new_n4159;
  assign new_n4215 = n2045 & new_n4153;
  assign new_n4216 = new_n4126 & new_n4215;
  assign new_n4217 = new_n4216 ^ new_n4214;
  assign new_n4218 = ~new_n4217 & new_n4123;
  assign new_n4219 = new_n4218 ^ new_n4217;
  assign new_n4220 = n2048 & new_n4153;
  assign new_n4221 = ~new_n4169 & new_n4220;
  assign new_n4222 = n2047 & new_n4153;
  assign new_n4223 = ~new_n4125 & ~new_n4222;
  assign new_n4224 = new_n4223 ^ new_n4169;
  assign new_n4225 = ~new_n4124 & ~new_n4222;
  assign new_n4226 = ~new_n4125 & ~new_n4225;
  assign new_n4227 = new_n4226 ^ new_n4224;
  assign new_n4228 = ~new_n4221 & new_n4227;
  assign new_n4229 = n2046 & new_n4153;
  assign new_n4230 = ~new_n4169 & new_n4229;
  assign new_n4231 = new_n4124 & new_n4220;
  assign new_n4232 = new_n4231 ^ new_n4124;
  assign new_n4233 = new_n4232 ^ new_n4220;
  assign new_n4234 = new_n4233 ^ new_n4124;
  assign new_n4235 = new_n4234 ^ new_n4230;
  assign new_n4236 = new_n4235 ^ new_n4228;
  assign new_n4237 = new_n4236 ^ new_n4123;
  assign new_n4238 = ~new_n4123 & ~new_n4236;
  assign new_n4239 = new_n4238 ^ new_n4237;
  assign new_n4240 = new_n4219 & new_n4239;
  assign new_n4241 = new_n4240 ^ new_n4122;
  assign new_n4242 = ~new_n4122 & new_n4240;
  assign new_n4243 = new_n4242 ^ new_n4241;
  assign new_n4244 = ~new_n4243 & new_n4207;
  assign new_n4245 = ~new_n4244 & new_n4121;
  assign new_n4246 = n2033 & new_n4152;
  assign new_n4247 = new_n4246 ^ new_n4121;
  assign new_n4248 = new_n4121 & new_n4246;
  assign new_n4249 = new_n4248 ^ new_n4247;
  assign new_n4250 = ~new_n4245 & new_n4249;
  assign new_n4251 = n2047 & new_n4118;
  assign new_n4252 = new_n4111 & new_n4251;
  assign new_n4253 = n2048 ^ n2047;
  assign new_n4254 = ~new_n4253 & new_n4118;
  assign new_n4255 = new_n4111 & new_n4254;
  assign new_n4256 = ~new_n4255 & new_n4252;
  assign new_n4257 = new_n4256 ^ new_n4252;
  assign new_n4258 = new_n4257 ^ new_n4255;
  assign new_n4259 = new_n4250 & new_n4258;
  assign new_n4260 = new_n4104 ^ new_n4098;
  assign new_n4261 = ~new_n4132 & new_n4260;
  assign new_n4262 = ~n2023 & ~n2024;
  assign new_n4263 = ~n2026 & ~n2027;
  assign new_n4264 = new_n4262 & new_n4263;
  assign new_n4265 = new_n4117 & new_n4264;
  assign new_n4266 = ~new_n4107 & new_n4265;
  assign new_n4267 = ~new_n4261 & ~new_n4266;
  assign new_n4268 = new_n4108 ^ n2044;
  assign new_n4269 = ~n2043 & ~new_n4268;
  assign new_n4270 = ~n2047 & new_n4269;
  assign new_n4271 = new_n4269 ^ new_n4268;
  assign new_n4272 = ~n2048 & n2046;
  assign new_n4273 = new_n4272 ^ n2048;
  assign new_n4274 = new_n4273 ^ new_n4113;
  assign new_n4275 = ~new_n4271 & ~new_n4274;
  assign new_n4276 = ~n2047 & n2048;
  assign new_n4277 = new_n4276 ^ new_n4272;
  assign new_n4278 = new_n4277 ^ new_n4114;
  assign new_n4279 = new_n4109 & new_n4278;
  assign new_n4280 = ~new_n4275 & ~new_n4279;
  assign new_n4281 = ~new_n4270 & new_n4280;
  assign new_n4282 = ~new_n4107 & ~new_n4281;
  assign new_n4283 = ~n2030 & ~n2031;
  assign new_n4284 = ~n2029 & new_n4283;
  assign new_n4285 = ~new_n4284 & new_n4106;
  assign new_n4286 = new_n4285 ^ new_n4106;
  assign new_n4287 = ~new_n4282 & ~new_n4286;
  assign new_n4288 = ~n2020 & new_n4287;
  assign new_n4289 = ~new_n4288 & new_n4118;
  assign new_n4290 = ~new_n4289 & new_n4267;
  assign new_n4291 = new_n4105 ^ n2021;
  assign new_n4292 = ~new_n4132 & ~new_n4291;
  assign new_n4293 = new_n4112 ^ n2046;
  assign new_n4294 = new_n4293 ^ new_n4274;
  assign new_n4295 = ~new_n4271 & new_n4294;
  assign new_n4296 = new_n4272 ^ n2047;
  assign new_n4297 = ~new_n4296 & new_n4109;
  assign new_n4298 = ~new_n4270 & ~new_n4297;
  assign new_n4299 = ~new_n4295 & new_n4298;
  assign new_n4300 = ~new_n4107 & ~new_n4299;
  assign new_n4301 = ~new_n4286 & ~new_n4300;
  assign new_n4302 = ~n2020 & new_n4301;
  assign new_n4303 = ~new_n4302 & new_n4118;
  assign new_n4304 = ~new_n4292 & ~new_n4303;
  assign new_n4305 = new_n4266 ^ new_n4151;
  assign new_n4306 = new_n4304 & new_n4305;
  assign new_n4307 = new_n4293 ^ new_n4272;
  assign new_n4308 = ~new_n4307 & new_n4109;
  assign new_n4309 = ~new_n4295 & ~new_n4308;
  assign new_n4310 = ~new_n4107 & ~new_n4309;
  assign new_n4311 = ~new_n4100 & ~new_n4310;
  assign new_n4312 = ~new_n4311 & new_n4118;
  assign new_n4313 = ~new_n4132 & new_n4105;
  assign new_n4314 = ~new_n4312 & ~new_n4313;
  assign new_n4315 = new_n4314 ^ new_n4306;
  assign new_n4316 = new_n4290 & new_n4315;
  assign new_n4317 = n2033 & new_n4153;
  assign new_n4318 = new_n4316 ^ new_n4315;
  assign new_n4319 = ~new_n4306 & ~new_n4314;
  assign new_n4320 = new_n4319 ^ new_n4314;
  assign new_n4321 = ~new_n4290 & ~new_n4320;
  assign new_n4322 = new_n4321 ^ new_n4318;
  assign new_n4323 = new_n4314 ^ new_n4290;
  assign new_n4324 = new_n4323 ^ new_n4322;
  assign new_n4325 = new_n4324 ^ new_n4317;
  assign new_n4326 = new_n4324 ^ new_n4196;
  assign new_n4327 = new_n4324 ^ new_n4193;
  assign new_n4328 = new_n4324 ^ new_n4187;
  assign new_n4329 = new_n4324 ^ new_n4184;
  assign new_n4330 = new_n4324 ^ new_n4175;
  assign new_n4331 = new_n4324 ^ new_n4172;
  assign new_n4332 = new_n4324 ^ new_n4162;
  assign new_n4333 = new_n4324 ^ new_n4155;
  assign new_n4334 = new_n4324 ^ new_n4157;
  assign new_n4335 = n2043 & new_n4153;
  assign new_n4336 = new_n4335 ^ new_n4324;
  assign new_n4337 = ~new_n4220 & ~new_n4324;
  assign new_n4338 = ~new_n4234 & ~new_n4337;
  assign new_n4339 = new_n4324 ^ new_n4222;
  assign new_n4340 = new_n4339 ^ new_n4338;
  assign new_n4341 = new_n4339 ^ new_n4125;
  assign new_n4342 = ~new_n4340 & new_n4341;
  assign new_n4343 = new_n4342 ^ new_n4125;
  assign new_n4344 = new_n4324 ^ new_n4229;
  assign new_n4345 = new_n4344 ^ new_n4343;
  assign new_n4346 = new_n4344 ^ new_n4123;
  assign new_n4347 = ~new_n4345 & new_n4346;
  assign new_n4348 = new_n4347 ^ new_n4123;
  assign new_n4349 = new_n4324 ^ new_n4215;
  assign new_n4350 = new_n4349 ^ new_n4348;
  assign new_n4351 = new_n4349 ^ new_n4122;
  assign new_n4352 = ~new_n4350 & new_n4351;
  assign new_n4353 = new_n4352 ^ new_n4122;
  assign new_n4354 = new_n4324 ^ new_n4208;
  assign new_n4355 = new_n4354 ^ new_n4353;
  assign new_n4356 = new_n4354 ^ new_n4121;
  assign new_n4357 = ~new_n4355 & new_n4356;
  assign new_n4358 = new_n4357 ^ new_n4121;
  assign new_n4359 = new_n4336 & new_n4358;
  assign new_n4360 = new_n4334 & new_n4359;
  assign new_n4361 = new_n4333 & new_n4360;
  assign new_n4362 = new_n4332 & new_n4361;
  assign new_n4363 = new_n4331 & new_n4362;
  assign new_n4364 = new_n4330 & new_n4363;
  assign new_n4365 = new_n4329 & new_n4364;
  assign new_n4366 = new_n4328 & new_n4365;
  assign new_n4367 = new_n4327 & new_n4366;
  assign new_n4368 = new_n4326 & new_n4367;
  assign new_n4369 = new_n4325 & new_n4368;
  assign new_n4370 = new_n4324 ^ new_n4246;
  assign new_n4371 = new_n4369 & new_n4370;
  assign new_n4372 = new_n4371 ^ new_n4370;
  assign new_n4373 = new_n4316 & new_n4372;
  assign new_n4374 = ~new_n4259 & ~new_n4373;
  assign new_n4375 = new_n4246 & new_n4257;
  assign new_n4376 = ~new_n4122 & new_n4121;
  assign new_n4377 = new_n4122 & new_n4123;
  assign new_n4378 = new_n4377 ^ new_n4123;
  assign new_n4379 = new_n4378 ^ new_n4376;
  assign new_n4380 = ~new_n4121 & new_n4378;
  assign new_n4381 = new_n4380 ^ new_n4379;
  assign new_n4382 = new_n4378 ^ new_n4122;
  assign new_n4383 = new_n4382 ^ new_n4381;
  assign new_n4384 = ~new_n4383 & new_n4256;
  assign new_n4385 = new_n4246 ^ new_n4125;
  assign new_n4386 = ~new_n4125 & ~new_n4246;
  assign new_n4387 = new_n4386 ^ new_n4385;
  assign new_n4388 = new_n4387 ^ new_n4246;
  assign new_n4389 = ~new_n4388 & new_n4384;
  assign new_n4390 = ~new_n4375 & ~new_n4389;
  assign new_n4391 = new_n4374 & new_n4390;
  assign new_n4392 = new_n4109 & new_n4251;
  assign new_n4393 = ~new_n4107 & n2046;
  assign new_n4394 = n2048 & new_n4393;
  assign new_n4395 = new_n4392 & new_n4394;
  assign new_n4396 = ~new_n4246 & new_n4395;
  assign new_n4397 = ~new_n4290 & new_n4319;
  assign new_n4398 = new_n4397 ^ new_n4322;
  assign new_n4399 = new_n4246 & new_n4398;
  assign new_n4400 = ~new_n4396 & ~new_n4399;
  assign new_n4401 = new_n4391 & new_n4400;
  assign new_n4402 = ~new_n4107 & ~new_n4270;
  assign new_n4403 = new_n4402 ^ new_n4147;
  assign new_n4404 = ~new_n4403 & new_n4118;
  assign new_n4405 = new_n4402 ^ new_n4285;
  assign new_n4406 = new_n4405 ^ new_n4098;
  assign new_n4407 = ~new_n4406 & new_n4118;
  assign new_n4408 = ~new_n4405 & new_n4118;
  assign new_n4409 = new_n4408 ^ new_n4407;
  assign new_n4410 = new_n4409 ^ new_n4404;
  assign new_n4411 = ~new_n4401 & new_n4410;
  assign new_n4412 = new_n4135 ^ new_n4107;
  assign new_n4413 = new_n4118 & new_n4412;
  assign new_n4414 = ~n2032 & new_n4284;
  assign new_n4415 = ~new_n4414 & new_n4106;
  assign new_n4416 = ~new_n4136 & ~new_n4415;
  assign new_n4417 = ~new_n4137 & new_n4416;
  assign new_n4418 = new_n4413 & new_n4417;
  assign new_n4419 = new_n4173 ^ new_n4163;
  assign new_n4420 = ~new_n4125 & new_n4419;
  assign new_n4421 = new_n4420 ^ new_n4419;
  assign new_n4422 = new_n4185 ^ new_n4176;
  assign new_n4423 = new_n4125 & new_n4422;
  assign new_n4424 = new_n4423 ^ new_n4422;
  assign new_n4425 = ~new_n4421 & ~new_n4424;
  assign new_n4426 = ~new_n4123 & ~new_n4425;
  assign new_n4427 = new_n4426 ^ new_n4425;
  assign new_n4428 = new_n4194 ^ new_n4188;
  assign new_n4429 = ~new_n4125 & new_n4428;
  assign new_n4430 = new_n4429 ^ new_n4428;
  assign new_n4431 = ~new_n4124 & ~new_n4317;
  assign new_n4432 = new_n4431 ^ new_n4197;
  assign new_n4433 = new_n4125 & new_n4432;
  assign new_n4434 = new_n4433 ^ new_n4432;
  assign new_n4435 = ~new_n4430 & ~new_n4434;
  assign new_n4436 = ~new_n4435 & new_n4123;
  assign new_n4437 = new_n4436 ^ new_n4435;
  assign new_n4438 = new_n4427 & new_n4437;
  assign new_n4439 = ~new_n4438 & new_n4122;
  assign new_n4440 = new_n4439 ^ new_n4438;
  assign new_n4441 = ~new_n4124 & ~new_n4335;
  assign new_n4442 = new_n4441 ^ new_n4211;
  assign new_n4443 = ~new_n4125 & new_n4442;
  assign new_n4444 = new_n4443 ^ new_n4442;
  assign new_n4445 = ~new_n4169 & new_n4155;
  assign new_n4446 = new_n4155 ^ new_n4125;
  assign new_n4447 = new_n4446 ^ new_n4445;
  assign new_n4448 = new_n4447 ^ new_n4154;
  assign new_n4449 = ~new_n4444 & new_n4448;
  assign new_n4450 = ~new_n4449 & new_n4123;
  assign new_n4451 = new_n4450 ^ new_n4449;
  assign new_n4452 = ~new_n4124 & ~new_n4215;
  assign new_n4453 = ~new_n4229 & new_n4124;
  assign new_n4454 = new_n4453 ^ new_n4452;
  assign new_n4455 = new_n4125 & new_n4454;
  assign new_n4456 = new_n4455 ^ new_n4454;
  assign new_n4457 = new_n4232 ^ new_n4225;
  assign new_n4458 = new_n4457 ^ new_n4125;
  assign new_n4459 = ~new_n4125 & ~new_n4457;
  assign new_n4460 = new_n4459 ^ new_n4458;
  assign new_n4461 = ~new_n4456 & new_n4460;
  assign new_n4462 = new_n4461 ^ new_n4123;
  assign new_n4463 = ~new_n4123 & new_n4461;
  assign new_n4464 = new_n4463 ^ new_n4462;
  assign new_n4465 = ~new_n4464 & new_n4451;
  assign new_n4466 = new_n4465 ^ new_n4122;
  assign new_n4467 = ~new_n4122 & new_n4465;
  assign new_n4468 = new_n4467 ^ new_n4466;
  assign new_n4469 = ~new_n4468 & new_n4440;
  assign new_n4470 = ~new_n4469 & new_n4121;
  assign new_n4471 = ~new_n4470 & new_n4249;
  assign new_n4472 = new_n4258 & new_n4471;
  assign new_n4473 = ~new_n4373 & ~new_n4472;
  assign new_n4474 = new_n4168 & new_n4246;
  assign new_n4475 = new_n4474 ^ new_n4388;
  assign new_n4476 = ~new_n4475 & new_n4384;
  assign new_n4477 = ~new_n4375 & ~new_n4476;
  assign new_n4478 = new_n4473 & new_n4477;
  assign new_n4479 = new_n4400 & new_n4478;
  assign new_n4480 = new_n4401 & new_n4479;
  assign new_n4481 = new_n4170 ^ new_n4125;
  assign new_n4482 = ~new_n4123 & ~new_n4481;
  assign new_n4483 = new_n4482 ^ new_n4481;
  assign new_n4484 = new_n4191 ^ new_n4179;
  assign new_n4485 = new_n4123 & new_n4484;
  assign new_n4486 = new_n4485 ^ new_n4484;
  assign new_n4487 = ~new_n4486 & new_n4483;
  assign new_n4488 = ~new_n4487 & new_n4122;
  assign new_n4489 = new_n4488 ^ new_n4487;
  assign new_n4490 = ~n2047 & new_n4124;
  assign new_n4491 = new_n4229 ^ new_n4157;
  assign new_n4492 = new_n4491 ^ new_n4159;
  assign new_n4493 = ~new_n4490 & new_n4492;
  assign new_n4494 = ~new_n4493 & new_n4125;
  assign new_n4495 = new_n4452 ^ new_n4215;
  assign new_n4496 = new_n4495 ^ new_n4212;
  assign new_n4497 = ~new_n4125 & new_n4496;
  assign new_n4498 = ~new_n4494 & ~new_n4497;
  assign new_n4499 = ~new_n4498 & new_n4123;
  assign new_n4500 = new_n4499 ^ new_n4498;
  assign new_n4501 = new_n4221 ^ new_n4123;
  assign new_n4502 = ~new_n4123 & new_n4221;
  assign new_n4503 = new_n4502 ^ new_n4501;
  assign new_n4504 = ~new_n4503 & new_n4500;
  assign new_n4505 = new_n4504 ^ new_n4122;
  assign new_n4506 = ~new_n4122 & new_n4504;
  assign new_n4507 = new_n4506 ^ new_n4505;
  assign new_n4508 = ~new_n4507 & new_n4489;
  assign new_n4509 = ~new_n4508 & new_n4121;
  assign new_n4510 = new_n4386 ^ new_n4200;
  assign new_n4511 = ~new_n4123 & new_n4510;
  assign new_n4512 = ~new_n4123 & ~new_n4246;
  assign new_n4513 = new_n4512 ^ new_n4510;
  assign new_n4514 = new_n4513 ^ new_n4511;
  assign new_n4515 = ~new_n4122 & new_n4514;
  assign new_n4516 = ~new_n4122 & new_n4246;
  assign new_n4517 = new_n4516 ^ new_n4122;
  assign new_n4518 = new_n4517 ^ new_n4514;
  assign new_n4519 = new_n4518 ^ new_n4515;
  assign new_n4520 = ~new_n4121 & ~new_n4519;
  assign new_n4521 = ~new_n4509 & ~new_n4520;
  assign new_n4522 = new_n4258 & new_n4521;
  assign new_n4523 = ~new_n4373 & ~new_n4522;
  assign new_n4524 = new_n4246 & new_n4384;
  assign new_n4525 = ~new_n4375 & ~new_n4524;
  assign new_n4526 = new_n4523 & new_n4525;
  assign new_n4527 = new_n4400 & new_n4526;
  assign new_n4528 = new_n4447 ^ new_n4420;
  assign new_n4529 = ~new_n4123 & new_n4528;
  assign new_n4530 = new_n4529 ^ new_n4528;
  assign new_n4531 = new_n4429 ^ new_n4423;
  assign new_n4532 = new_n4123 & new_n4531;
  assign new_n4533 = new_n4532 ^ new_n4531;
  assign new_n4534 = ~new_n4530 & ~new_n4533;
  assign new_n4535 = ~new_n4534 & new_n4122;
  assign new_n4536 = new_n4535 ^ new_n4534;
  assign new_n4537 = new_n4455 ^ new_n4443;
  assign new_n4538 = new_n4123 & new_n4537;
  assign new_n4539 = new_n4538 ^ new_n4537;
  assign new_n4540 = new_n4459 ^ new_n4123;
  assign new_n4541 = ~new_n4123 & new_n4459;
  assign new_n4542 = new_n4541 ^ new_n4540;
  assign new_n4543 = ~new_n4539 & ~new_n4542;
  assign new_n4544 = new_n4543 ^ new_n4122;
  assign new_n4545 = ~new_n4122 & new_n4543;
  assign new_n4546 = new_n4545 ^ new_n4544;
  assign new_n4547 = ~new_n4546 & new_n4536;
  assign new_n4548 = ~new_n4547 & new_n4121;
  assign new_n4549 = new_n4433 ^ new_n4386;
  assign new_n4550 = ~new_n4123 & new_n4549;
  assign new_n4551 = new_n4549 ^ new_n4512;
  assign new_n4552 = new_n4551 ^ new_n4550;
  assign new_n4553 = ~new_n4122 & new_n4552;
  assign new_n4554 = new_n4552 ^ new_n4517;
  assign new_n4555 = new_n4554 ^ new_n4553;
  assign new_n4556 = ~new_n4121 & ~new_n4555;
  assign new_n4557 = ~new_n4548 & ~new_n4556;
  assign new_n4558 = new_n4258 & new_n4557;
  assign new_n4559 = ~new_n4373 & ~new_n4558;
  assign new_n4560 = new_n4126 & new_n4246;
  assign new_n4561 = new_n4560 ^ new_n4246;
  assign new_n4562 = new_n4384 & new_n4561;
  assign new_n4563 = ~new_n4375 & ~new_n4562;
  assign new_n4564 = new_n4559 & new_n4563;
  assign new_n4565 = new_n4400 & new_n4564;
  assign new_n4566 = new_n4527 & new_n4565;
  assign new_n4567 = new_n4480 & new_n4566;
  assign new_n4568 = new_n4218 ^ new_n4182;
  assign new_n4569 = new_n4122 & new_n4568;
  assign new_n4570 = new_n4238 ^ new_n4122;
  assign new_n4571 = ~new_n4122 & new_n4238;
  assign new_n4572 = new_n4571 ^ new_n4570;
  assign new_n4573 = new_n4572 ^ new_n4568;
  assign new_n4574 = new_n4573 ^ new_n4569;
  assign new_n4575 = new_n4121 & new_n4574;
  assign new_n4576 = new_n4512 ^ new_n4203;
  assign new_n4577 = ~new_n4122 & new_n4576;
  assign new_n4578 = new_n4576 ^ new_n4517;
  assign new_n4579 = new_n4578 ^ new_n4577;
  assign new_n4580 = ~new_n4121 & ~new_n4579;
  assign new_n4581 = ~new_n4575 & ~new_n4580;
  assign new_n4582 = new_n4258 & new_n4581;
  assign new_n4583 = ~new_n4373 & ~new_n4582;
  assign new_n4584 = ~new_n4388 & new_n4378;
  assign new_n4585 = ~new_n4377 & new_n4246;
  assign new_n4586 = new_n4585 ^ new_n4516;
  assign new_n4587 = new_n4512 ^ new_n4123;
  assign new_n4588 = new_n4587 ^ new_n4586;
  assign new_n4589 = ~new_n4584 & new_n4588;
  assign new_n4590 = ~new_n4589 & new_n4121;
  assign new_n4591 = new_n4590 ^ new_n4589;
  assign new_n4592 = ~new_n4591 & new_n4256;
  assign new_n4593 = ~new_n4375 & ~new_n4592;
  assign new_n4594 = new_n4583 & new_n4593;
  assign new_n4595 = new_n4400 & new_n4594;
  assign new_n4596 = new_n4450 ^ new_n4426;
  assign new_n4597 = new_n4122 & new_n4596;
  assign new_n4598 = new_n4597 ^ new_n4596;
  assign new_n4599 = ~new_n4122 & new_n4463;
  assign new_n4600 = new_n4599 ^ new_n4122;
  assign new_n4601 = new_n4600 ^ new_n4463;
  assign new_n4602 = ~new_n4598 & ~new_n4601;
  assign new_n4603 = ~new_n4602 & new_n4121;
  assign new_n4604 = new_n4512 ^ new_n4436;
  assign new_n4605 = ~new_n4122 & new_n4604;
  assign new_n4606 = new_n4604 ^ new_n4517;
  assign new_n4607 = new_n4606 ^ new_n4605;
  assign new_n4608 = ~new_n4121 & ~new_n4607;
  assign new_n4609 = ~new_n4603 & ~new_n4608;
  assign new_n4610 = new_n4258 & new_n4609;
  assign new_n4611 = ~new_n4373 & ~new_n4610;
  assign new_n4612 = new_n4475 & new_n4587;
  assign new_n4613 = ~new_n4612 & new_n4256;
  assign new_n4614 = new_n4122 ^ new_n4121;
  assign new_n4615 = new_n4614 ^ new_n4376;
  assign new_n4616 = new_n4615 ^ new_n4121;
  assign new_n4617 = ~new_n4616 & new_n4613;
  assign new_n4618 = ~new_n4375 & ~new_n4617;
  assign new_n4619 = new_n4611 & new_n4618;
  assign new_n4620 = new_n4400 & new_n4619;
  assign new_n4621 = new_n4595 & new_n4620;
  assign new_n4622 = new_n4502 ^ new_n4122;
  assign new_n4623 = ~new_n4122 & new_n4502;
  assign new_n4624 = new_n4623 ^ new_n4622;
  assign new_n4625 = new_n4499 ^ new_n4482;
  assign new_n4626 = new_n4625 ^ new_n4624;
  assign new_n4627 = new_n4122 & new_n4625;
  assign new_n4628 = new_n4627 ^ new_n4626;
  assign new_n4629 = new_n4121 & new_n4628;
  assign new_n4630 = new_n4511 ^ new_n4485;
  assign new_n4631 = ~new_n4122 & new_n4630;
  assign new_n4632 = new_n4630 ^ new_n4517;
  assign new_n4633 = new_n4632 ^ new_n4631;
  assign new_n4634 = ~new_n4121 & ~new_n4633;
  assign new_n4635 = ~new_n4629 & ~new_n4634;
  assign new_n4636 = new_n4258 & new_n4635;
  assign new_n4637 = ~new_n4373 & ~new_n4636;
  assign new_n4638 = new_n4121 & new_n4516;
  assign new_n4639 = new_n4638 ^ new_n4516;
  assign new_n4640 = new_n4256 & new_n4639;
  assign new_n4641 = ~new_n4375 & ~new_n4640;
  assign new_n4642 = new_n4637 & new_n4641;
  assign new_n4643 = new_n4400 & new_n4642;
  assign new_n4644 = new_n4538 ^ new_n4529;
  assign new_n4645 = new_n4122 & new_n4644;
  assign new_n4646 = new_n4645 ^ new_n4644;
  assign new_n4647 = new_n4541 ^ new_n4122;
  assign new_n4648 = ~new_n4122 & new_n4541;
  assign new_n4649 = new_n4648 ^ new_n4647;
  assign new_n4650 = ~new_n4646 & ~new_n4649;
  assign new_n4651 = ~new_n4650 & new_n4121;
  assign new_n4652 = new_n4550 ^ new_n4532;
  assign new_n4653 = ~new_n4122 & new_n4652;
  assign new_n4654 = new_n4652 ^ new_n4517;
  assign new_n4655 = new_n4654 ^ new_n4653;
  assign new_n4656 = ~new_n4121 & ~new_n4655;
  assign new_n4657 = ~new_n4651 & ~new_n4656;
  assign new_n4658 = new_n4258 & new_n4657;
  assign new_n4659 = ~new_n4373 & ~new_n4658;
  assign new_n4660 = new_n4378 & new_n4561;
  assign new_n4661 = ~new_n4660 & new_n4588;
  assign new_n4662 = ~new_n4661 & new_n4121;
  assign new_n4663 = new_n4662 ^ new_n4661;
  assign new_n4664 = ~new_n4663 & new_n4256;
  assign new_n4665 = ~new_n4375 & ~new_n4664;
  assign new_n4666 = new_n4659 & new_n4665;
  assign new_n4667 = new_n4400 & new_n4666;
  assign new_n4668 = new_n4643 & new_n4667;
  assign new_n4669 = new_n4621 & new_n4668;
  assign new_n4670 = new_n4567 & new_n4669;
  assign new_n4671 = ~new_n4242 & new_n4121;
  assign new_n4672 = new_n4517 ^ new_n4206;
  assign new_n4673 = ~new_n4121 & ~new_n4672;
  assign new_n4674 = ~new_n4671 & ~new_n4673;
  assign new_n4675 = new_n4258 & new_n4674;
  assign new_n4676 = ~new_n4373 & ~new_n4675;
  assign new_n4677 = new_n4377 ^ new_n4122;
  assign new_n4678 = ~new_n4388 & new_n4677;
  assign new_n4679 = ~new_n4516 & ~new_n4678;
  assign new_n4680 = ~new_n4679 & new_n4121;
  assign new_n4681 = new_n4680 ^ new_n4679;
  assign new_n4682 = ~new_n4681 & new_n4256;
  assign new_n4683 = ~new_n4375 & ~new_n4682;
  assign new_n4684 = new_n4676 & new_n4683;
  assign new_n4685 = new_n4400 & new_n4684;
  assign new_n4686 = ~new_n4467 & new_n4121;
  assign new_n4687 = new_n4517 ^ new_n4439;
  assign new_n4688 = ~new_n4121 & ~new_n4687;
  assign new_n4689 = ~new_n4686 & ~new_n4688;
  assign new_n4690 = new_n4258 & new_n4689;
  assign new_n4691 = ~new_n4373 & ~new_n4690;
  assign new_n4692 = ~new_n4475 & new_n4677;
  assign new_n4693 = ~new_n4516 & ~new_n4692;
  assign new_n4694 = ~new_n4693 & new_n4121;
  assign new_n4695 = new_n4694 ^ new_n4693;
  assign new_n4696 = ~new_n4695 & new_n4256;
  assign new_n4697 = ~new_n4375 & ~new_n4696;
  assign new_n4698 = new_n4691 & new_n4697;
  assign new_n4699 = new_n4400 & new_n4698;
  assign new_n4700 = new_n4685 & new_n4699;
  assign new_n4701 = ~new_n4506 & new_n4121;
  assign new_n4702 = new_n4515 ^ new_n4488;
  assign new_n4703 = ~new_n4121 & new_n4702;
  assign new_n4704 = ~new_n4701 & ~new_n4703;
  assign new_n4705 = new_n4258 & new_n4704;
  assign new_n4706 = ~new_n4373 & ~new_n4705;
  assign new_n4707 = ~new_n4123 & new_n4615;
  assign new_n4708 = new_n4246 & new_n4707;
  assign new_n4709 = new_n4249 ^ new_n4121;
  assign new_n4710 = new_n4709 ^ new_n4708;
  assign new_n4711 = new_n4710 ^ new_n4639;
  assign new_n4712 = new_n4711 ^ new_n4248;
  assign new_n4713 = new_n4712 ^ new_n4246;
  assign new_n4714 = new_n4256 & new_n4713;
  assign new_n4715 = ~new_n4375 & ~new_n4714;
  assign new_n4716 = new_n4706 & new_n4715;
  assign new_n4717 = new_n4400 & new_n4716;
  assign new_n4718 = ~new_n4545 & new_n4121;
  assign new_n4719 = new_n4553 ^ new_n4535;
  assign new_n4720 = ~new_n4121 & new_n4719;
  assign new_n4721 = ~new_n4718 & ~new_n4720;
  assign new_n4722 = new_n4258 & new_n4721;
  assign new_n4723 = ~new_n4373 & ~new_n4722;
  assign new_n4724 = new_n4561 & new_n4677;
  assign new_n4725 = ~new_n4516 & ~new_n4724;
  assign new_n4726 = ~new_n4725 & new_n4121;
  assign new_n4727 = new_n4726 ^ new_n4725;
  assign new_n4728 = ~new_n4727 & new_n4256;
  assign new_n4729 = ~new_n4375 & ~new_n4728;
  assign new_n4730 = new_n4723 & new_n4729;
  assign new_n4731 = new_n4400 & new_n4730;
  assign new_n4732 = new_n4717 & new_n4731;
  assign new_n4733 = new_n4700 & new_n4732;
  assign new_n4734 = ~new_n4571 & new_n4121;
  assign new_n4735 = new_n4577 ^ new_n4569;
  assign new_n4736 = ~new_n4121 & new_n4735;
  assign new_n4737 = ~new_n4734 & ~new_n4736;
  assign new_n4738 = new_n4258 & new_n4737;
  assign new_n4739 = ~new_n4373 & ~new_n4738;
  assign new_n4740 = ~new_n4585 & new_n4475;
  assign new_n4741 = ~new_n4474 & new_n4740;
  assign new_n4742 = ~new_n4741 & new_n4121;
  assign new_n4743 = new_n4742 ^ new_n4741;
  assign new_n4744 = ~new_n4743 & new_n4256;
  assign new_n4745 = ~new_n4375 & ~new_n4744;
  assign new_n4746 = new_n4739 & new_n4745;
  assign new_n4747 = new_n4400 & new_n4746;
  assign new_n4748 = ~new_n4599 & new_n4121;
  assign new_n4749 = new_n4605 ^ new_n4597;
  assign new_n4750 = ~new_n4121 & new_n4749;
  assign new_n4751 = ~new_n4748 & ~new_n4750;
  assign new_n4752 = new_n4258 & new_n4751;
  assign new_n4753 = ~new_n4373 & ~new_n4752;
  assign new_n4754 = ~new_n4740 & new_n4121;
  assign new_n4755 = new_n4754 ^ new_n4740;
  assign new_n4756 = ~new_n4755 & new_n4256;
  assign new_n4757 = ~new_n4375 & ~new_n4756;
  assign new_n4758 = new_n4753 & new_n4757;
  assign new_n4759 = new_n4400 & new_n4758;
  assign new_n4760 = new_n4747 & new_n4759;
  assign new_n4761 = new_n4370 ^ new_n4369;
  assign new_n4762 = new_n4316 & new_n4761;
  assign new_n4763 = ~new_n4623 & new_n4121;
  assign new_n4764 = new_n4631 ^ new_n4627;
  assign new_n4765 = ~new_n4121 & new_n4764;
  assign new_n4766 = ~new_n4763 & ~new_n4765;
  assign new_n4767 = new_n4258 & new_n4766;
  assign new_n4768 = ~new_n4762 & ~new_n4767;
  assign new_n4769 = new_n4256 & new_n4709;
  assign new_n4770 = ~new_n4375 & ~new_n4769;
  assign new_n4771 = new_n4768 & new_n4770;
  assign new_n4772 = new_n4400 & new_n4771;
  assign new_n4773 = ~new_n4648 & new_n4121;
  assign new_n4774 = new_n4653 ^ new_n4645;
  assign new_n4775 = ~new_n4121 & new_n4774;
  assign new_n4776 = ~new_n4773 & ~new_n4775;
  assign new_n4777 = new_n4258 & new_n4776;
  assign new_n4778 = ~new_n4373 & ~new_n4777;
  assign new_n4779 = ~new_n4561 & ~new_n4585;
  assign new_n4780 = ~new_n4779 & new_n4121;
  assign new_n4781 = new_n4780 ^ new_n4779;
  assign new_n4782 = ~new_n4781 & new_n4256;
  assign new_n4783 = ~new_n4375 & ~new_n4782;
  assign new_n4784 = new_n4778 & new_n4783;
  assign new_n4785 = new_n4400 & new_n4784;
  assign new_n4786 = new_n4772 & new_n4785;
  assign new_n4787 = new_n4760 & new_n4786;
  assign new_n4788 = new_n4733 & new_n4787;
  assign new_n4789 = new_n4670 & new_n4788;
  assign new_n4790 = new_n4367 ^ new_n4326;
  assign new_n4791 = new_n4316 & new_n4790;
  assign new_n4792 = ~new_n4121 & new_n4258;
  assign new_n4793 = new_n4244 & new_n4792;
  assign new_n4794 = ~new_n4791 & ~new_n4793;
  assign new_n4795 = ~new_n4388 & new_n4381;
  assign new_n4796 = ~new_n4711 & ~new_n4795;
  assign new_n4797 = new_n4168 & new_n4317;
  assign new_n4798 = new_n4126 ^ new_n4125;
  assign new_n4799 = new_n4196 & new_n4798;
  assign new_n4800 = new_n4799 ^ new_n4124;
  assign new_n4801 = new_n4800 ^ new_n4198;
  assign new_n4802 = ~new_n4797 & ~new_n4801;
  assign new_n4803 = new_n4387 & new_n4802;
  assign new_n4804 = ~new_n4383 & ~new_n4803;
  assign new_n4805 = new_n4246 & new_n4381;
  assign new_n4806 = new_n4805 ^ new_n4588;
  assign new_n4807 = new_n4806 ^ new_n4713;
  assign new_n4808 = ~new_n4804 & new_n4807;
  assign new_n4809 = new_n4796 & new_n4808;
  assign new_n4810 = ~new_n4809 & new_n4256;
  assign new_n4811 = new_n4808 ^ new_n4712;
  assign new_n4812 = ~new_n4811 & new_n4257;
  assign new_n4813 = ~new_n4810 & ~new_n4812;
  assign new_n4814 = new_n4794 & new_n4813;
  assign new_n4815 = ~new_n4196 & new_n4395;
  assign new_n4816 = new_n4196 & new_n4398;
  assign new_n4817 = ~new_n4815 & ~new_n4816;
  assign new_n4818 = new_n4814 & new_n4817;
  assign new_n4819 = new_n4368 ^ new_n4325;
  assign new_n4820 = new_n4316 & new_n4819;
  assign new_n4821 = new_n4469 & new_n4792;
  assign new_n4822 = ~new_n4820 & ~new_n4821;
  assign new_n4823 = ~new_n4475 & new_n4381;
  assign new_n4824 = ~new_n4711 & ~new_n4823;
  assign new_n4825 = new_n4317 & new_n4798;
  assign new_n4826 = new_n4825 ^ new_n4124;
  assign new_n4827 = new_n4826 ^ new_n4431;
  assign new_n4828 = ~new_n4474 & new_n4827;
  assign new_n4829 = new_n4387 & new_n4828;
  assign new_n4830 = ~new_n4383 & ~new_n4829;
  assign new_n4831 = new_n4830 ^ new_n4807;
  assign new_n4832 = new_n4824 & new_n4831;
  assign new_n4833 = ~new_n4832 & new_n4256;
  assign new_n4834 = new_n4830 ^ new_n4712;
  assign new_n4835 = ~new_n4834 & new_n4807;
  assign new_n4836 = ~new_n4835 & new_n4257;
  assign new_n4837 = ~new_n4833 & ~new_n4836;
  assign new_n4838 = new_n4822 & new_n4837;
  assign new_n4839 = ~new_n4317 & new_n4395;
  assign new_n4840 = new_n4317 & new_n4398;
  assign new_n4841 = ~new_n4839 & ~new_n4840;
  assign new_n4842 = new_n4838 & new_n4841;
  assign new_n4843 = new_n4818 & new_n4842;
  assign new_n4844 = new_n4365 ^ new_n4328;
  assign new_n4845 = new_n4316 & new_n4844;
  assign new_n4846 = new_n4508 & new_n4792;
  assign new_n4847 = ~new_n4845 & ~new_n4846;
  assign new_n4848 = new_n4126 & new_n4317;
  assign new_n4849 = ~new_n4799 & ~new_n4848;
  assign new_n4850 = new_n4195 ^ new_n4189;
  assign new_n4851 = ~new_n4850 & new_n4125;
  assign new_n4852 = new_n4851 ^ new_n4850;
  assign new_n4853 = new_n4849 & new_n4852;
  assign new_n4854 = ~new_n4383 & ~new_n4853;
  assign new_n4855 = ~new_n4854 & new_n4807;
  assign new_n4856 = new_n4805 ^ new_n4711;
  assign new_n4857 = ~new_n4856 & new_n4855;
  assign new_n4858 = ~new_n4857 & new_n4256;
  assign new_n4859 = new_n4855 ^ new_n4712;
  assign new_n4860 = ~new_n4859 & new_n4257;
  assign new_n4861 = ~new_n4858 & ~new_n4860;
  assign new_n4862 = new_n4847 & new_n4861;
  assign new_n4863 = ~new_n4187 & new_n4395;
  assign new_n4864 = new_n4187 & new_n4398;
  assign new_n4865 = ~new_n4863 & ~new_n4864;
  assign new_n4866 = new_n4862 & new_n4865;
  assign new_n4867 = new_n4366 ^ new_n4327;
  assign new_n4868 = new_n4316 & new_n4867;
  assign new_n4869 = new_n4547 & new_n4792;
  assign new_n4870 = ~new_n4868 & ~new_n4869;
  assign new_n4871 = new_n4381 & new_n4561;
  assign new_n4872 = ~new_n4711 & ~new_n4871;
  assign new_n4873 = new_n4197 ^ new_n4194;
  assign new_n4874 = ~new_n4873 & new_n4125;
  assign new_n4875 = new_n4874 ^ new_n4873;
  assign new_n4876 = new_n4825 ^ new_n4560;
  assign new_n4877 = ~new_n4876 & new_n4875;
  assign new_n4878 = ~new_n4383 & ~new_n4877;
  assign new_n4879 = ~new_n4878 & new_n4807;
  assign new_n4880 = new_n4872 & new_n4879;
  assign new_n4881 = ~new_n4880 & new_n4256;
  assign new_n4882 = new_n4879 ^ new_n4712;
  assign new_n4883 = ~new_n4882 & new_n4257;
  assign new_n4884 = ~new_n4881 & ~new_n4883;
  assign new_n4885 = new_n4870 & new_n4884;
  assign new_n4886 = ~new_n4193 & new_n4395;
  assign new_n4887 = new_n4193 & new_n4398;
  assign new_n4888 = ~new_n4886 & ~new_n4887;
  assign new_n4889 = new_n4885 & new_n4888;
  assign new_n4890 = new_n4866 & new_n4889;
  assign new_n4891 = new_n4843 & new_n4890;
  assign new_n4892 = new_n4363 ^ new_n4330;
  assign new_n4893 = new_n4316 & new_n4892;
  assign new_n4894 = ~new_n4574 & new_n4792;
  assign new_n4895 = ~new_n4893 & ~new_n4894;
  assign new_n4896 = ~new_n4803 & new_n4380;
  assign new_n4897 = ~new_n4708 & ~new_n4896;
  assign new_n4898 = new_n4186 ^ new_n4177;
  assign new_n4899 = new_n4898 ^ new_n4851;
  assign new_n4900 = ~new_n4898 & new_n4125;
  assign new_n4901 = new_n4900 ^ new_n4899;
  assign new_n4902 = ~new_n4383 & ~new_n4901;
  assign new_n4903 = ~new_n4590 & ~new_n4902;
  assign new_n4904 = ~new_n4711 & new_n4903;
  assign new_n4905 = new_n4897 & new_n4904;
  assign new_n4906 = ~new_n4905 & new_n4256;
  assign new_n4907 = ~new_n4712 & ~new_n4902;
  assign new_n4908 = new_n4897 & new_n4907;
  assign new_n4909 = ~new_n4908 & new_n4257;
  assign new_n4910 = ~new_n4906 & ~new_n4909;
  assign new_n4911 = new_n4895 & new_n4910;
  assign new_n4912 = ~new_n4175 & new_n4395;
  assign new_n4913 = new_n4175 & new_n4398;
  assign new_n4914 = ~new_n4912 & ~new_n4913;
  assign new_n4915 = new_n4911 & new_n4914;
  assign new_n4916 = new_n4364 ^ new_n4329;
  assign new_n4917 = new_n4316 & new_n4916;
  assign new_n4918 = new_n4602 & new_n4792;
  assign new_n4919 = ~new_n4917 & ~new_n4918;
  assign new_n4920 = ~new_n4612 & new_n4376;
  assign new_n4921 = ~new_n4711 & ~new_n4920;
  assign new_n4922 = new_n4188 ^ new_n4185;
  assign new_n4923 = new_n4922 ^ new_n4874;
  assign new_n4924 = ~new_n4922 & new_n4125;
  assign new_n4925 = new_n4924 ^ new_n4923;
  assign new_n4926 = ~new_n4383 & ~new_n4925;
  assign new_n4927 = ~new_n4829 & new_n4380;
  assign new_n4928 = ~new_n4708 & ~new_n4927;
  assign new_n4929 = ~new_n4926 & new_n4928;
  assign new_n4930 = new_n4921 & new_n4929;
  assign new_n4931 = ~new_n4930 & new_n4256;
  assign new_n4932 = new_n4929 ^ new_n4712;
  assign new_n4933 = ~new_n4932 & new_n4257;
  assign new_n4934 = ~new_n4931 & ~new_n4933;
  assign new_n4935 = new_n4919 & new_n4934;
  assign new_n4936 = ~new_n4184 & new_n4395;
  assign new_n4937 = new_n4184 & new_n4398;
  assign new_n4938 = ~new_n4936 & ~new_n4937;
  assign new_n4939 = new_n4935 & new_n4938;
  assign new_n4940 = new_n4915 & new_n4939;
  assign new_n4941 = new_n4361 ^ new_n4332;
  assign new_n4942 = new_n4316 & new_n4941;
  assign new_n4943 = ~new_n4628 & new_n4792;
  assign new_n4944 = ~new_n4942 & ~new_n4943;
  assign new_n4945 = ~new_n4853 & new_n4380;
  assign new_n4946 = ~new_n4708 & ~new_n4945;
  assign new_n4947 = new_n4166 & new_n4174;
  assign new_n4948 = new_n4174 ^ new_n4164;
  assign new_n4949 = new_n4948 ^ new_n4947;
  assign new_n4950 = ~new_n4900 & new_n4949;
  assign new_n4951 = ~new_n4383 & ~new_n4950;
  assign new_n4952 = new_n4951 ^ new_n4638;
  assign new_n4953 = ~new_n4711 & ~new_n4952;
  assign new_n4954 = new_n4946 & new_n4953;
  assign new_n4955 = ~new_n4954 & new_n4256;
  assign new_n4956 = new_n4946 ^ new_n4712;
  assign new_n4957 = new_n4956 ^ new_n4951;
  assign new_n4958 = ~new_n4957 & new_n4257;
  assign new_n4959 = ~new_n4955 & ~new_n4958;
  assign new_n4960 = new_n4944 & new_n4959;
  assign new_n4961 = ~new_n4162 & new_n4395;
  assign new_n4962 = new_n4162 & new_n4398;
  assign new_n4963 = ~new_n4961 & ~new_n4962;
  assign new_n4964 = new_n4960 & new_n4963;
  assign new_n4965 = new_n4362 ^ new_n4331;
  assign new_n4966 = new_n4316 & new_n4965;
  assign new_n4967 = new_n4650 & new_n4792;
  assign new_n4968 = ~new_n4966 & ~new_n4967;
  assign new_n4969 = ~new_n4877 & new_n4380;
  assign new_n4970 = ~new_n4708 & ~new_n4969;
  assign new_n4971 = new_n4176 ^ new_n4173;
  assign new_n4972 = new_n4971 ^ new_n4924;
  assign new_n4973 = ~new_n4971 & new_n4125;
  assign new_n4974 = new_n4973 ^ new_n4972;
  assign new_n4975 = ~new_n4383 & ~new_n4974;
  assign new_n4976 = ~new_n4662 & ~new_n4975;
  assign new_n4977 = ~new_n4711 & new_n4976;
  assign new_n4978 = new_n4970 & new_n4977;
  assign new_n4979 = ~new_n4978 & new_n4256;
  assign new_n4980 = ~new_n4712 & ~new_n4975;
  assign new_n4981 = new_n4970 & new_n4980;
  assign new_n4982 = ~new_n4981 & new_n4257;
  assign new_n4983 = ~new_n4979 & ~new_n4982;
  assign new_n4984 = new_n4968 & new_n4983;
  assign new_n4985 = ~new_n4172 & new_n4395;
  assign new_n4986 = new_n4172 & new_n4398;
  assign new_n4987 = ~new_n4985 & ~new_n4986;
  assign new_n4988 = new_n4984 & new_n4987;
  assign new_n4989 = new_n4964 & new_n4988;
  assign new_n4990 = new_n4940 & new_n4989;
  assign new_n4991 = new_n4891 & new_n4990;
  assign new_n4992 = new_n4359 ^ new_n4334;
  assign new_n4993 = new_n4316 & new_n4992;
  assign new_n4994 = new_n4242 & new_n4792;
  assign new_n4995 = ~new_n4993 & ~new_n4994;
  assign new_n4996 = ~new_n4901 & new_n4380;
  assign new_n4997 = ~new_n4803 & new_n4707;
  assign new_n4998 = ~new_n4996 & ~new_n4997;
  assign new_n4999 = new_n4680 ^ new_n4159;
  assign new_n5000 = new_n4999 ^ new_n4711;
  assign new_n5001 = ~new_n5000 & new_n4998;
  assign new_n5002 = ~new_n5001 & new_n4256;
  assign new_n5003 = ~new_n4159 & ~new_n4712;
  assign new_n5004 = new_n4998 & new_n5003;
  assign new_n5005 = ~new_n5004 & new_n4257;
  assign new_n5006 = ~new_n5002 & ~new_n5005;
  assign new_n5007 = new_n4995 & new_n5006;
  assign new_n5008 = ~new_n4157 & new_n4395;
  assign new_n5009 = new_n4157 & new_n4398;
  assign new_n5010 = ~new_n5008 & ~new_n5009;
  assign new_n5011 = new_n5007 & new_n5010;
  assign new_n5012 = new_n4360 ^ new_n4333;
  assign new_n5013 = new_n4316 & new_n5012;
  assign new_n5014 = new_n4467 & new_n4792;
  assign new_n5015 = ~new_n5013 & ~new_n5014;
  assign new_n5016 = ~new_n4925 & new_n4380;
  assign new_n5017 = ~new_n4829 & new_n4707;
  assign new_n5018 = ~new_n5016 & ~new_n5017;
  assign new_n5019 = new_n4694 ^ new_n4445;
  assign new_n5020 = ~new_n4711 & ~new_n5019;
  assign new_n5021 = new_n5018 & new_n5020;
  assign new_n5022 = ~new_n5021 & new_n4256;
  assign new_n5023 = ~new_n4445 & ~new_n4712;
  assign new_n5024 = new_n5018 & new_n5023;
  assign new_n5025 = ~new_n5024 & new_n4257;
  assign new_n5026 = ~new_n5022 & ~new_n5025;
  assign new_n5027 = new_n5015 & new_n5026;
  assign new_n5028 = ~new_n4155 & new_n4395;
  assign new_n5029 = new_n4155 & new_n4398;
  assign new_n5030 = ~new_n5028 & ~new_n5029;
  assign new_n5031 = new_n5027 & new_n5030;
  assign new_n5032 = new_n5011 & new_n5031;
  assign new_n5033 = new_n4222 ^ new_n4125;
  assign new_n5034 = new_n5033 ^ new_n4223;
  assign new_n5035 = ~new_n5034 & new_n4321;
  assign new_n5036 = new_n4397 & new_n5033;
  assign new_n5037 = ~new_n5035 & ~new_n5036;
  assign new_n5038 = ~new_n4223 & new_n4322;
  assign new_n5039 = new_n4223 & new_n4395;
  assign new_n5040 = ~new_n5038 & ~new_n5039;
  assign new_n5041 = new_n5037 & new_n5040;
  assign new_n5042 = new_n4340 ^ new_n4125;
  assign new_n5043 = new_n4316 & new_n5042;
  assign new_n5044 = new_n4648 & new_n4792;
  assign new_n5045 = ~new_n5043 & ~new_n5044;
  assign new_n5046 = new_n4707 ^ new_n4615;
  assign new_n5047 = ~new_n4877 & new_n5046;
  assign new_n5048 = ~new_n4453 & new_n4226;
  assign new_n5049 = ~new_n4125 & ~new_n4452;
  assign new_n5050 = ~new_n4211 & new_n5049;
  assign new_n5051 = new_n4452 ^ new_n4211;
  assign new_n5052 = new_n5051 ^ new_n5050;
  assign new_n5053 = ~new_n5048 & new_n5052;
  assign new_n5054 = ~new_n4383 & ~new_n5053;
  assign new_n5055 = ~new_n5047 & ~new_n5054;
  assign new_n5056 = ~new_n4974 & new_n4707;
  assign new_n5057 = new_n4126 & new_n4162;
  assign new_n5058 = new_n4160 ^ new_n4155;
  assign new_n5059 = new_n5058 ^ new_n4445;
  assign new_n5060 = ~new_n5057 & ~new_n5059;
  assign new_n5061 = new_n4335 & new_n4798;
  assign new_n5062 = new_n5061 ^ new_n4124;
  assign new_n5063 = new_n5062 ^ new_n4441;
  assign new_n5064 = ~new_n4156 & new_n5063;
  assign new_n5065 = new_n5060 & new_n5064;
  assign new_n5066 = ~new_n5065 & new_n4380;
  assign new_n5067 = new_n5066 ^ new_n4780;
  assign new_n5068 = ~new_n5056 & ~new_n5067;
  assign new_n5069 = new_n5055 & new_n5068;
  assign new_n5070 = ~new_n5069 & new_n4256;
  assign new_n5071 = new_n5066 ^ new_n4248;
  assign new_n5072 = ~new_n5056 & ~new_n5071;
  assign new_n5073 = new_n5055 & new_n5072;
  assign new_n5074 = ~new_n5073 & new_n4257;
  assign new_n5075 = ~new_n5070 & ~new_n5074;
  assign new_n5076 = new_n5045 & new_n5075;
  assign new_n5077 = new_n5041 & new_n5076;
  assign new_n5078 = new_n4220 ^ new_n4124;
  assign new_n5079 = new_n4397 & new_n5078;
  assign new_n5080 = new_n4233 & new_n4322;
  assign new_n5081 = ~new_n4233 & new_n4395;
  assign new_n5082 = ~new_n5080 & ~new_n5081;
  assign new_n5083 = ~new_n5079 & new_n5082;
  assign new_n5084 = new_n4231 & new_n4321;
  assign new_n5085 = new_n4316 & new_n5078;
  assign new_n5086 = ~new_n5084 & ~new_n5085;
  assign new_n5087 = new_n5083 & new_n5086;
  assign new_n5088 = ~new_n4246 & new_n4372;
  assign new_n5089 = new_n4321 ^ new_n4290;
  assign new_n5090 = new_n5089 ^ new_n4398;
  assign new_n5091 = ~new_n5090 & new_n5088;
  assign new_n5092 = new_n4397 ^ new_n4319;
  assign new_n5093 = ~new_n4371 & new_n5092;
  assign new_n5094 = ~new_n5091 & ~new_n5093;
  assign new_n5095 = new_n4623 & new_n4792;
  assign new_n5096 = ~new_n4853 & new_n5046;
  assign new_n5097 = new_n4229 & new_n4798;
  assign new_n5098 = ~new_n4216 & ~new_n5097;
  assign new_n5099 = new_n4228 & new_n5098;
  assign new_n5100 = ~new_n4383 & ~new_n5099;
  assign new_n5101 = ~new_n5096 & ~new_n5100;
  assign new_n5102 = new_n4168 & new_n4335;
  assign new_n5103 = ~new_n4209 & ~new_n5102;
  assign new_n5104 = ~new_n4160 & new_n5103;
  assign new_n5105 = ~new_n5104 & new_n4380;
  assign new_n5106 = ~new_n4248 & ~new_n5105;
  assign new_n5107 = ~new_n4950 & new_n4707;
  assign new_n5108 = ~new_n5107 & new_n5106;
  assign new_n5109 = new_n5101 & new_n5108;
  assign new_n5110 = ~new_n5109 & new_n4252;
  assign new_n5111 = ~new_n5095 & ~new_n5110;
  assign new_n5112 = new_n5094 & new_n5111;
  assign new_n5113 = new_n5087 & new_n5112;
  assign new_n5114 = ~new_n5077 & ~new_n5113;
  assign new_n5115 = new_n5114 ^ new_n5113;
  assign new_n5116 = new_n5115 ^ new_n5077;
  assign new_n5117 = ~new_n5116 & new_n5032;
  assign new_n5118 = new_n4358 ^ new_n4336;
  assign new_n5119 = new_n4316 & new_n5118;
  assign new_n5120 = new_n4545 & new_n4792;
  assign new_n5121 = ~new_n5119 & ~new_n5120;
  assign new_n5122 = ~new_n4974 & new_n4380;
  assign new_n5123 = ~new_n4877 & new_n4707;
  assign new_n5124 = ~new_n5122 & ~new_n5123;
  assign new_n5125 = ~new_n4383 & ~new_n5065;
  assign new_n5126 = ~new_n4726 & ~new_n5125;
  assign new_n5127 = ~new_n4711 & new_n5126;
  assign new_n5128 = new_n5124 & new_n5127;
  assign new_n5129 = ~new_n5128 & new_n4256;
  assign new_n5130 = ~new_n4248 & ~new_n5125;
  assign new_n5131 = ~new_n4711 & new_n5130;
  assign new_n5132 = new_n5124 & new_n5131;
  assign new_n5133 = ~new_n5132 & new_n4257;
  assign new_n5134 = ~new_n5129 & ~new_n5133;
  assign new_n5135 = new_n5121 & new_n5134;
  assign new_n5136 = ~new_n4335 & new_n4395;
  assign new_n5137 = new_n4335 & new_n4398;
  assign new_n5138 = ~new_n5136 & ~new_n5137;
  assign new_n5139 = new_n5135 & new_n5138;
  assign new_n5140 = ~new_n4121 & ~new_n4208;
  assign new_n5141 = ~new_n5140 & new_n4322;
  assign new_n5142 = new_n4395 & new_n5140;
  assign new_n5143 = ~new_n5141 & ~new_n5142;
  assign new_n5144 = new_n4208 ^ new_n4121;
  assign new_n5145 = new_n4397 & new_n5144;
  assign new_n5146 = ~new_n5145 & new_n5143;
  assign new_n5147 = new_n4258 & new_n4506;
  assign new_n5148 = ~new_n4121 & ~new_n5147;
  assign new_n5149 = new_n4208 & new_n4321;
  assign new_n5150 = ~new_n5149 & new_n4121;
  assign new_n5151 = ~new_n5148 & ~new_n5150;
  assign new_n5152 = ~new_n5151 & new_n5146;
  assign new_n5153 = ~new_n4950 & new_n4380;
  assign new_n5154 = ~new_n4853 & new_n4707;
  assign new_n5155 = ~new_n5153 & ~new_n5154;
  assign new_n5156 = ~new_n4383 & ~new_n5104;
  assign new_n5157 = new_n4713 ^ new_n4585;
  assign new_n5158 = ~new_n5156 & ~new_n5157;
  assign new_n5159 = ~new_n4711 & new_n5158;
  assign new_n5160 = new_n5155 & new_n5159;
  assign new_n5161 = ~new_n5160 & new_n4256;
  assign new_n5162 = ~new_n4248 & ~new_n5156;
  assign new_n5163 = ~new_n4711 & new_n5162;
  assign new_n5164 = new_n5155 & new_n5163;
  assign new_n5165 = ~new_n5164 & new_n4257;
  assign new_n5166 = ~new_n5161 & ~new_n5165;
  assign new_n5167 = new_n4355 ^ new_n4121;
  assign new_n5168 = new_n4316 & new_n5167;
  assign new_n5169 = ~new_n5168 & new_n5166;
  assign new_n5170 = new_n5152 & new_n5169;
  assign new_n5171 = ~new_n4123 & ~new_n4229;
  assign new_n5172 = new_n4229 ^ new_n4123;
  assign new_n5173 = new_n5172 ^ new_n5171;
  assign new_n5174 = ~new_n5173 & new_n4321;
  assign new_n5175 = new_n4397 & new_n5172;
  assign new_n5176 = ~new_n5174 & ~new_n5175;
  assign new_n5177 = ~new_n5171 & new_n4322;
  assign new_n5178 = new_n4395 & new_n5171;
  assign new_n5179 = ~new_n5177 & ~new_n5178;
  assign new_n5180 = new_n5176 & new_n5179;
  assign new_n5181 = new_n4345 ^ new_n4123;
  assign new_n5182 = new_n4316 & new_n5181;
  assign new_n5183 = new_n4571 & new_n4792;
  assign new_n5184 = ~new_n5182 & ~new_n5183;
  assign new_n5185 = ~new_n4803 & new_n5046;
  assign new_n5186 = new_n4126 & new_n4335;
  assign new_n5187 = ~new_n4213 & ~new_n5186;
  assign new_n5188 = new_n4216 ^ new_n4124;
  assign new_n5189 = new_n5188 ^ new_n4495;
  assign new_n5190 = new_n5189 ^ new_n4230;
  assign new_n5191 = new_n5187 & new_n5190;
  assign new_n5192 = ~new_n4383 & ~new_n5191;
  assign new_n5193 = ~new_n5185 & ~new_n5192;
  assign new_n5194 = ~new_n4901 & new_n4707;
  assign new_n5195 = new_n4947 ^ new_n4159;
  assign new_n5196 = new_n4380 & new_n5195;
  assign new_n5197 = new_n5196 ^ new_n4742;
  assign new_n5198 = ~new_n5194 & ~new_n5197;
  assign new_n5199 = new_n5193 & new_n5198;
  assign new_n5200 = ~new_n5199 & new_n4256;
  assign new_n5201 = new_n5196 ^ new_n4248;
  assign new_n5202 = ~new_n5194 & ~new_n5201;
  assign new_n5203 = new_n5193 & new_n5202;
  assign new_n5204 = ~new_n5203 & new_n4257;
  assign new_n5205 = ~new_n5200 & ~new_n5204;
  assign new_n5206 = new_n5184 & new_n5205;
  assign new_n5207 = new_n5180 & new_n5206;
  assign new_n5208 = ~new_n4122 & ~new_n4215;
  assign new_n5209 = new_n4215 ^ new_n4122;
  assign new_n5210 = new_n5209 ^ new_n5208;
  assign new_n5211 = ~new_n5210 & new_n4321;
  assign new_n5212 = new_n4397 & new_n5209;
  assign new_n5213 = ~new_n5211 & ~new_n5212;
  assign new_n5214 = ~new_n5208 & new_n4322;
  assign new_n5215 = new_n4395 & new_n5208;
  assign new_n5216 = ~new_n5214 & ~new_n5215;
  assign new_n5217 = new_n5213 & new_n5216;
  assign new_n5218 = new_n4350 ^ new_n4122;
  assign new_n5219 = new_n4316 & new_n5218;
  assign new_n5220 = new_n4599 & new_n4792;
  assign new_n5221 = ~new_n5219 & ~new_n5220;
  assign new_n5222 = ~new_n4829 & new_n5046;
  assign new_n5223 = new_n5061 ^ new_n5050;
  assign new_n5224 = new_n5223 ^ new_n4160;
  assign new_n5225 = ~new_n4383 & new_n5224;
  assign new_n5226 = ~new_n5222 & ~new_n5225;
  assign new_n5227 = ~new_n4925 & new_n4707;
  assign new_n5228 = new_n5057 ^ new_n4124;
  assign new_n5229 = new_n5228 ^ new_n4163;
  assign new_n5230 = ~new_n4445 & ~new_n5229;
  assign new_n5231 = ~new_n4973 & new_n5230;
  assign new_n5232 = ~new_n5231 & new_n4380;
  assign new_n5233 = new_n5232 ^ new_n4754;
  assign new_n5234 = ~new_n5227 & ~new_n5233;
  assign new_n5235 = new_n5226 & new_n5234;
  assign new_n5236 = ~new_n5235 & new_n4256;
  assign new_n5237 = new_n5232 ^ new_n4248;
  assign new_n5238 = ~new_n5227 & ~new_n5237;
  assign new_n5239 = new_n5226 & new_n5238;
  assign new_n5240 = ~new_n5239 & new_n4257;
  assign new_n5241 = ~new_n5236 & ~new_n5240;
  assign new_n5242 = new_n5221 & new_n5241;
  assign new_n5243 = new_n5217 & new_n5242;
  assign new_n5244 = new_n5207 & new_n5243;
  assign new_n5245 = ~new_n5170 & new_n5244;
  assign new_n5246 = new_n5245 ^ new_n5244;
  assign new_n5247 = new_n5139 & new_n5246;
  assign new_n5248 = new_n5117 & new_n5247;
  assign new_n5249 = new_n4991 & new_n5248;
  assign new_n5250 = new_n4789 & new_n5249;
  assign new_n5251 = new_n4101 ^ n2020;
  assign new_n5252 = ~new_n5251 & new_n4408;
  assign new_n5253 = ~new_n5250 & ~new_n5252;
  assign new_n5254 = ~new_n5253 & new_n4418;
  assign new_n5255 = new_n4136 ^ new_n4100;
  assign new_n5256 = ~new_n5255 & new_n4413;
  assign new_n5257 = new_n5252 ^ new_n4418;
  assign new_n5258 = new_n4418 & new_n5252;
  assign new_n5259 = new_n5258 ^ new_n5257;
  assign new_n5260 = ~new_n5256 & new_n5259;
  assign new_n5261 = ~new_n5254 & new_n5260;
  assign new_n5262 = ~new_n4418 & new_n5256;
  assign new_n5263 = new_n4479 & new_n5262;
  assign new_n5264 = ~new_n5263 & new_n5252;
  assign new_n5265 = new_n5262 ^ new_n5256;
  assign new_n5266 = new_n5250 & new_n5265;
  assign new_n5267 = ~new_n5252 & ~new_n5266;
  assign new_n5268 = ~new_n5264 & ~new_n5267;
  assign new_n5269 = ~new_n5261 & ~new_n5268;
  assign new_n5270 = ~new_n4479 & new_n5265;
  assign new_n5271 = new_n5250 & new_n5258;
  assign new_n5272 = ~new_n5263 & ~new_n5271;
  assign new_n5273 = new_n5250 & new_n5256;
  assign new_n5274 = ~new_n5272 & ~new_n5273;
  assign new_n5275 = ~new_n5270 & ~new_n5274;
  assign new_n5276 = new_n5269 & new_n5275;
  assign new_n5277 = ~new_n5276 & n2033;
  assign new_n5278 = new_n4408 ^ new_n4404;
  assign new_n5279 = new_n5277 & new_n5278;
  assign new_n5280 = ~new_n4411 & ~new_n5279;
  assign new_n5281 = ~new_n4565 & new_n4410;
  assign new_n5282 = ~new_n5279 & ~new_n5281;
  assign new_n5283 = ~new_n4527 & new_n4410;
  assign new_n5284 = ~new_n5279 & ~new_n5283;
  assign new_n5285 = ~new_n4620 & new_n4410;
  assign new_n5286 = ~new_n5279 & ~new_n5285;
  assign new_n5287 = n2023 & new_n4409;
  assign new_n5288 = ~new_n5287 & new_n5286;
  assign new_n5289 = ~new_n4595 & new_n4410;
  assign new_n5290 = ~new_n5279 & ~new_n5289;
  assign new_n5291 = n2024 & new_n4409;
  assign new_n5292 = ~new_n5291 & new_n5290;
  assign new_n5293 = ~new_n4667 & new_n4410;
  assign new_n5294 = ~new_n5279 & ~new_n5293;
  assign new_n5295 = n2025 & new_n4409;
  assign new_n5296 = ~new_n5295 & new_n5294;
  assign new_n5297 = ~new_n4643 & new_n4410;
  assign new_n5298 = ~new_n5279 & ~new_n5297;
  assign new_n5299 = n2026 & new_n4409;
  assign new_n5300 = ~new_n5299 & new_n5298;
  assign new_n5301 = ~new_n4699 & new_n4410;
  assign new_n5302 = ~new_n5279 & ~new_n5301;
  assign new_n5303 = n2027 & new_n4409;
  assign new_n5304 = ~new_n5303 & new_n5302;
  assign new_n5305 = ~new_n4685 & new_n4410;
  assign new_n5306 = ~new_n5279 & ~new_n5305;
  assign new_n5307 = n2028 & new_n4409;
  assign new_n5308 = ~new_n5307 & new_n5306;
  assign new_n5309 = ~new_n4731 & new_n4410;
  assign new_n5310 = ~new_n5279 & ~new_n5309;
  assign new_n5311 = n2029 & new_n4409;
  assign new_n5312 = ~new_n5311 & new_n5310;
  assign new_n5313 = ~new_n4717 & new_n4410;
  assign new_n5314 = ~new_n5279 & ~new_n5313;
  assign new_n5315 = n2030 & new_n4409;
  assign new_n5316 = ~new_n5315 & new_n5314;
  assign new_n5317 = ~new_n4759 & new_n4410;
  assign new_n5318 = ~new_n5279 & ~new_n5317;
  assign new_n5319 = n2031 & new_n4409;
  assign new_n5320 = ~new_n5319 & new_n5318;
  assign new_n5321 = ~new_n4747 & new_n4410;
  assign new_n5322 = ~new_n5279 & ~new_n5321;
  assign new_n5323 = n2032 & new_n4409;
  assign new_n5324 = ~new_n5323 & new_n5322;
  assign new_n5325 = ~new_n4785 & new_n4410;
  assign new_n5326 = ~new_n5279 & ~new_n5325;
  assign new_n5327 = n2033 & new_n4409;
  assign new_n5328 = ~new_n5327 & new_n5326;
  assign new_n5329 = ~new_n4772 & new_n4410;
  assign new_n5330 = n2034 & new_n5278;
  assign new_n5331 = ~new_n5276 & new_n5330;
  assign new_n5332 = ~new_n5329 & ~new_n5331;
  assign new_n5333 = n2034 & new_n4409;
  assign new_n5334 = ~new_n5333 & new_n5332;
  assign new_n5335 = ~new_n4842 & new_n4410;
  assign new_n5336 = n2035 & new_n5278;
  assign new_n5337 = ~new_n5276 & new_n5336;
  assign new_n5338 = ~new_n5335 & ~new_n5337;
  assign new_n5339 = n2035 & new_n4409;
  assign new_n5340 = ~new_n5339 & new_n5338;
  assign new_n5341 = ~new_n4818 & new_n4410;
  assign new_n5342 = n2036 & new_n5278;
  assign new_n5343 = ~new_n5276 & new_n5342;
  assign new_n5344 = ~new_n5341 & ~new_n5343;
  assign new_n5345 = n2036 & new_n4409;
  assign new_n5346 = ~new_n5345 & new_n5344;
  assign new_n5347 = ~new_n4889 & new_n4410;
  assign new_n5348 = n2037 & new_n5278;
  assign new_n5349 = ~new_n5276 & new_n5348;
  assign new_n5350 = ~new_n5347 & ~new_n5349;
  assign new_n5351 = n2037 & new_n4409;
  assign new_n5352 = ~new_n5351 & new_n5350;
  assign new_n5353 = ~new_n4866 & new_n4410;
  assign new_n5354 = n2038 & new_n5278;
  assign new_n5355 = ~new_n5276 & new_n5354;
  assign new_n5356 = ~new_n5353 & ~new_n5355;
  assign new_n5357 = n2038 & new_n4409;
  assign new_n5358 = ~new_n5357 & new_n5356;
  assign new_n5359 = ~new_n4939 & new_n4410;
  assign new_n5360 = n2039 & new_n5278;
  assign new_n5361 = ~new_n5276 & new_n5360;
  assign new_n5362 = ~new_n5359 & ~new_n5361;
  assign new_n5363 = n2039 & new_n4409;
  assign new_n5364 = ~new_n5363 & new_n5362;
  assign new_n5365 = ~new_n4915 & new_n4410;
  assign new_n5366 = n2040 & new_n5278;
  assign new_n5367 = ~new_n5276 & new_n5366;
  assign new_n5368 = ~new_n5365 & ~new_n5367;
  assign new_n5369 = n2040 & new_n4409;
  assign new_n5370 = ~new_n5369 & new_n5368;
  assign new_n5371 = ~new_n4988 & new_n4410;
  assign new_n5372 = n2041 & new_n5278;
  assign new_n5373 = ~new_n5276 & new_n5372;
  assign new_n5374 = ~new_n5371 & ~new_n5373;
  assign new_n5375 = n2041 & new_n4409;
  assign new_n5376 = ~new_n5375 & new_n5374;
  assign new_n5377 = ~new_n4964 & new_n4410;
  assign new_n5378 = n2042 & new_n5278;
  assign new_n5379 = ~new_n5276 & new_n5378;
  assign new_n5380 = ~new_n5377 & ~new_n5379;
  assign new_n5381 = n2042 & new_n4409;
  assign new_n5382 = ~new_n5381 & new_n5380;
  assign new_n5383 = ~new_n5031 & new_n4410;
  assign new_n5384 = n2043 & new_n5278;
  assign new_n5385 = ~new_n5276 & new_n5384;
  assign new_n5386 = ~new_n5383 & ~new_n5385;
  assign new_n5387 = n2043 & new_n4409;
  assign new_n5388 = ~new_n5387 & new_n5386;
  assign new_n5389 = ~new_n5011 & new_n4410;
  assign new_n5390 = n2044 & new_n5278;
  assign new_n5391 = ~new_n5276 & new_n5390;
  assign new_n5392 = ~new_n5389 & ~new_n5391;
  assign new_n5393 = n2044 & new_n4409;
  assign new_n5394 = ~new_n5393 & new_n5392;
  assign new_n5395 = ~new_n5139 & new_n4410;
  assign new_n5396 = n2045 & new_n5278;
  assign new_n5397 = ~new_n5276 & new_n5396;
  assign new_n5398 = ~new_n5395 & ~new_n5397;
  assign new_n5399 = n2045 & new_n4409;
  assign new_n5400 = ~new_n5399 & new_n5398;
  assign new_n5401 = ~new_n5170 & new_n4410;
  assign new_n5402 = n2046 & new_n5278;
  assign new_n5403 = ~new_n5276 & new_n5402;
  assign new_n5404 = ~new_n5401 & ~new_n5403;
  assign new_n5405 = n2046 & new_n4409;
  assign new_n5406 = ~new_n5405 & new_n5404;
  assign new_n5407 = ~new_n5243 & new_n4410;
  assign new_n5408 = n2047 & new_n5278;
  assign new_n5409 = ~new_n5276 & new_n5408;
  assign new_n5410 = ~new_n5407 & ~new_n5409;
  assign new_n5411 = n2047 & new_n4409;
  assign new_n5412 = ~new_n5411 & new_n5410;
  assign new_n5413 = ~new_n4479 & new_n4410;
  assign new_n5414 = ~new_n5279 & ~new_n5413;
  assign new_n5415 = ~new_n5207 & new_n4410;
  assign new_n5416 = ~n2048 & ~new_n5276;
  assign new_n5417 = ~new_n5416 & new_n5278;
  assign new_n5418 = ~new_n5415 & ~new_n5417;
  assign new_n5419 = ~n2048 & new_n4404;
  assign new_n5420 = ~new_n4407 & ~new_n5419;
  assign new_n5421 = ~new_n5420 & new_n5418;
  assign new_n5422 = ~new_n5207 & ~new_n5243;
  assign new_n5423 = new_n5170 & new_n5422;
  assign new_n5424 = new_n5423 ^ new_n5422;
  assign new_n5425 = ~new_n5011 & ~new_n5139;
  assign new_n5426 = new_n5031 & new_n5425;
  assign new_n5427 = new_n5426 ^ new_n5425;
  assign new_n5428 = new_n5424 & new_n5427;
  assign new_n5429 = ~n2020 & new_n4140;
  assign new_n5430 = new_n5429 ^ new_n4141;
  assign new_n5431 = new_n5428 & new_n5430;
  assign new_n5432 = new_n5429 ^ new_n4148;
  assign new_n5433 = ~new_n5077 & new_n5432;
  assign new_n5434 = new_n5433 ^ new_n5432;
  assign new_n5435 = new_n5428 & new_n5434;
  assign new_n5436 = ~new_n5431 & ~new_n5435;
  assign new_n5437 = new_n5432 ^ new_n4141;
  assign new_n5438 = ~new_n5116 & new_n5437;
  assign new_n5439 = new_n5428 & new_n5438;
  assign new_n5440 = ~new_n5439 & new_n5436;
  assign new_n5441 = n2080 & new_n5440;
  assign new_n5442 = n2079 & new_n5440;
  assign new_n5443 = n2078 & new_n5440;
  assign new_n5444 = n2077 & new_n5440;
  assign new_n5445 = n2076 & new_n5440;
  assign new_n5446 = n2075 & new_n5440;
  assign new_n5447 = n2074 & new_n5440;
  assign new_n5448 = n2073 & new_n5440;
  assign new_n5449 = new_n5428 & new_n5437;
  assign new_n5450 = ~new_n5115 & new_n5449;
  assign new_n5451 = ~new_n5450 & new_n5436;
  assign new_n5452 = n2072 & new_n5451;
  assign new_n5453 = n2071 & new_n5451;
  assign new_n5454 = n2070 & new_n5451;
  assign new_n5455 = n2069 & new_n5451;
  assign new_n5456 = n2068 & new_n5451;
  assign new_n5457 = n2067 & new_n5451;
  assign new_n5458 = n2066 & new_n5451;
  assign new_n5459 = n2065 & new_n5451;
  assign new_n5460 = new_n5428 & new_n5433;
  assign new_n5461 = ~new_n5431 & ~new_n5460;
  assign new_n5462 = new_n5114 ^ new_n5077;
  assign new_n5463 = ~new_n5462 & new_n5449;
  assign new_n5464 = ~new_n5463 & new_n5461;
  assign new_n5465 = n2064 & new_n5464;
  assign new_n5466 = n2063 & new_n5464;
  assign new_n5467 = n2062 & new_n5464;
  assign new_n5468 = n2061 & new_n5464;
  assign new_n5469 = n2060 & new_n5464;
  assign new_n5470 = n2059 & new_n5464;
  assign new_n5471 = n2058 & new_n5464;
  assign new_n5472 = n2057 & new_n5464;
  assign new_n5473 = new_n5114 & new_n5449;
  assign new_n5474 = ~new_n5473 & new_n5461;
  assign new_n5475 = n2056 & new_n5474;
  assign new_n5476 = n2055 & new_n5474;
  assign new_n5477 = n2054 & new_n5474;
  assign new_n5478 = n2053 & new_n5474;
  assign new_n5479 = n2052 & new_n5474;
  assign new_n5480 = n2051 & new_n5474;
  assign new_n5481 = n2050 & new_n5474;
  assign new_n5482 = n2049 & new_n5474;
  assign new_n5483 = ~new_n5243 & new_n5207;
  assign new_n5484 = new_n5170 & new_n5483;
  assign new_n5485 = new_n5484 ^ new_n5483;
  assign new_n5486 = new_n5427 & new_n5485;
  assign new_n5487 = new_n5430 & new_n5486;
  assign new_n5488 = new_n5434 & new_n5486;
  assign new_n5489 = ~new_n5487 & ~new_n5488;
  assign new_n5490 = new_n5438 & new_n5486;
  assign new_n5491 = ~new_n5490 & new_n5489;
  assign new_n5492 = n2112 & new_n5491;
  assign new_n5493 = n2111 & new_n5491;
  assign new_n5494 = n2110 & new_n5491;
  assign new_n5495 = n2109 & new_n5491;
  assign new_n5496 = n2108 & new_n5491;
  assign new_n5497 = n2107 & new_n5491;
  assign new_n5498 = n2106 & new_n5491;
  assign new_n5499 = n2105 & new_n5491;
  assign new_n5500 = ~new_n5115 & new_n5437;
  assign new_n5501 = new_n5486 & new_n5500;
  assign new_n5502 = ~new_n5501 & new_n5489;
  assign new_n5503 = n2104 & new_n5502;
  assign new_n5504 = n2103 & new_n5502;
  assign new_n5505 = n2102 & new_n5502;
  assign new_n5506 = n2101 & new_n5502;
  assign new_n5507 = n2100 & new_n5502;
  assign new_n5508 = n2099 & new_n5502;
  assign new_n5509 = n2098 & new_n5502;
  assign new_n5510 = n2097 & new_n5502;
  assign new_n5511 = new_n5433 & new_n5486;
  assign new_n5512 = ~new_n5487 & ~new_n5511;
  assign new_n5513 = ~new_n5462 & new_n5437;
  assign new_n5514 = new_n5486 & new_n5513;
  assign new_n5515 = ~new_n5514 & new_n5512;
  assign new_n5516 = n2096 & new_n5515;
  assign new_n5517 = n2095 & new_n5515;
  assign new_n5518 = n2094 & new_n5515;
  assign new_n5519 = n2093 & new_n5515;
  assign new_n5520 = n2092 & new_n5515;
  assign new_n5521 = n2091 & new_n5515;
  assign new_n5522 = n2090 & new_n5515;
  assign new_n5523 = n2089 & new_n5515;
  assign new_n5524 = new_n5114 & new_n5437;
  assign new_n5525 = new_n5486 & new_n5524;
  assign new_n5526 = ~new_n5525 & new_n5512;
  assign new_n5527 = n2088 & new_n5526;
  assign new_n5528 = n2087 & new_n5526;
  assign new_n5529 = n2086 & new_n5526;
  assign new_n5530 = n2085 & new_n5526;
  assign new_n5531 = n2084 & new_n5526;
  assign new_n5532 = n2083 & new_n5526;
  assign new_n5533 = n2082 & new_n5526;
  assign new_n5534 = n2081 & new_n5526;
  assign new_n5535 = ~new_n5207 & new_n5243;
  assign new_n5536 = new_n5170 & new_n5535;
  assign new_n5537 = new_n5536 ^ new_n5535;
  assign new_n5538 = new_n5427 & new_n5537;
  assign new_n5539 = new_n5434 & new_n5538;
  assign new_n5540 = new_n5430 & new_n5538;
  assign new_n5541 = ~new_n5539 & ~new_n5540;
  assign new_n5542 = new_n5438 & new_n5538;
  assign new_n5543 = ~new_n5542 & new_n5541;
  assign new_n5544 = n2144 & new_n5543;
  assign new_n5545 = n2143 & new_n5543;
  assign new_n5546 = n2142 & new_n5543;
  assign new_n5547 = n2141 & new_n5543;
  assign new_n5548 = n2140 & new_n5543;
  assign new_n5549 = n2139 & new_n5543;
  assign new_n5550 = n2138 & new_n5543;
  assign new_n5551 = n2137 & new_n5543;
  assign new_n5552 = new_n5500 & new_n5538;
  assign new_n5553 = ~new_n5552 & new_n5541;
  assign new_n5554 = n2136 & new_n5553;
  assign new_n5555 = n2135 & new_n5553;
  assign new_n5556 = n2134 & new_n5553;
  assign new_n5557 = n2133 & new_n5553;
  assign new_n5558 = n2132 & new_n5553;
  assign new_n5559 = n2131 & new_n5553;
  assign new_n5560 = n2130 & new_n5553;
  assign new_n5561 = n2129 & new_n5553;
  assign new_n5562 = new_n5433 & new_n5538;
  assign new_n5563 = ~new_n5540 & ~new_n5562;
  assign new_n5564 = new_n5513 & new_n5538;
  assign new_n5565 = ~new_n5564 & new_n5563;
  assign new_n5566 = n2128 & new_n5565;
  assign new_n5567 = n2127 & new_n5565;
  assign new_n5568 = n2126 & new_n5565;
  assign new_n5569 = n2125 & new_n5565;
  assign new_n5570 = n2124 & new_n5565;
  assign new_n5571 = n2123 & new_n5565;
  assign new_n5572 = n2122 & new_n5565;
  assign new_n5573 = n2121 & new_n5565;
  assign new_n5574 = new_n5524 & new_n5538;
  assign new_n5575 = ~new_n5574 & new_n5563;
  assign new_n5576 = n2120 & new_n5575;
  assign new_n5577 = n2119 & new_n5575;
  assign new_n5578 = n2118 & new_n5575;
  assign new_n5579 = n2117 & new_n5575;
  assign new_n5580 = n2116 & new_n5575;
  assign new_n5581 = n2115 & new_n5575;
  assign new_n5582 = n2114 & new_n5575;
  assign new_n5583 = n2113 & new_n5575;
  assign new_n5584 = new_n5245 & new_n5427;
  assign new_n5585 = new_n5434 & new_n5584;
  assign new_n5586 = new_n5430 & new_n5584;
  assign new_n5587 = ~new_n5585 & ~new_n5586;
  assign new_n5588 = new_n5438 & new_n5584;
  assign new_n5589 = ~new_n5588 & new_n5587;
  assign new_n5590 = n2176 & new_n5589;
  assign new_n5591 = n2175 & new_n5589;
  assign new_n5592 = n2174 & new_n5589;
  assign new_n5593 = n2173 & new_n5589;
  assign new_n5594 = n2172 & new_n5589;
  assign new_n5595 = n2171 & new_n5589;
  assign new_n5596 = n2170 & new_n5589;
  assign new_n5597 = n2169 & new_n5589;
  assign new_n5598 = new_n5500 & new_n5584;
  assign new_n5599 = ~new_n5598 & new_n5587;
  assign new_n5600 = n2168 & new_n5599;
  assign new_n5601 = n2167 & new_n5599;
  assign new_n5602 = n2166 & new_n5599;
  assign new_n5603 = n2165 & new_n5599;
  assign new_n5604 = n2164 & new_n5599;
  assign new_n5605 = n2163 & new_n5599;
  assign new_n5606 = n2162 & new_n5599;
  assign new_n5607 = n2161 & new_n5599;
  assign new_n5608 = new_n5433 & new_n5584;
  assign new_n5609 = ~new_n5586 & ~new_n5608;
  assign new_n5610 = new_n5513 & new_n5584;
  assign new_n5611 = ~new_n5610 & new_n5609;
  assign new_n5612 = n2160 & new_n5611;
  assign new_n5613 = n2159 & new_n5611;
  assign new_n5614 = n2158 & new_n5611;
  assign new_n5615 = n2157 & new_n5611;
  assign new_n5616 = n2156 & new_n5611;
  assign new_n5617 = n2155 & new_n5611;
  assign new_n5618 = n2154 & new_n5611;
  assign new_n5619 = n2153 & new_n5611;
  assign new_n5620 = new_n5524 & new_n5584;
  assign new_n5621 = ~new_n5620 & new_n5609;
  assign new_n5622 = n2152 & new_n5621;
  assign new_n5623 = n2151 & new_n5621;
  assign new_n5624 = n2150 & new_n5621;
  assign new_n5625 = n2149 & new_n5621;
  assign new_n5626 = n2148 & new_n5621;
  assign new_n5627 = n2147 & new_n5621;
  assign new_n5628 = n2146 & new_n5621;
  assign new_n5629 = n2145 & new_n5621;
  assign new_n5630 = new_n5423 & new_n5427;
  assign new_n5631 = new_n5434 & new_n5630;
  assign new_n5632 = new_n5430 & new_n5630;
  assign new_n5633 = ~new_n5631 & ~new_n5632;
  assign new_n5634 = new_n5438 & new_n5630;
  assign new_n5635 = ~new_n5634 & new_n5633;
  assign new_n5636 = n2208 & new_n5635;
  assign new_n5637 = n2207 & new_n5635;
  assign new_n5638 = n2206 & new_n5635;
  assign new_n5639 = n2205 & new_n5635;
  assign new_n5640 = n2204 & new_n5635;
  assign new_n5641 = n2203 & new_n5635;
  assign new_n5642 = n2202 & new_n5635;
  assign new_n5643 = n2201 & new_n5635;
  assign new_n5644 = new_n5500 & new_n5630;
  assign new_n5645 = ~new_n5644 & new_n5633;
  assign new_n5646 = n2200 & new_n5645;
  assign new_n5647 = n2199 & new_n5645;
  assign new_n5648 = n2198 & new_n5645;
  assign new_n5649 = n2197 & new_n5645;
  assign new_n5650 = n2196 & new_n5645;
  assign new_n5651 = n2195 & new_n5645;
  assign new_n5652 = n2194 & new_n5645;
  assign new_n5653 = n2193 & new_n5645;
  assign new_n5654 = new_n5433 & new_n5630;
  assign new_n5655 = ~new_n5632 & ~new_n5654;
  assign new_n5656 = new_n5513 & new_n5630;
  assign new_n5657 = ~new_n5656 & new_n5655;
  assign new_n5658 = n2192 & new_n5657;
  assign new_n5659 = n2191 & new_n5657;
  assign new_n5660 = n2190 & new_n5657;
  assign new_n5661 = n2189 & new_n5657;
  assign new_n5662 = n2188 & new_n5657;
  assign new_n5663 = n2187 & new_n5657;
  assign new_n5664 = n2186 & new_n5657;
  assign new_n5665 = n2185 & new_n5657;
  assign new_n5666 = new_n5524 & new_n5630;
  assign new_n5667 = ~new_n5666 & new_n5655;
  assign new_n5668 = n2184 & new_n5667;
  assign new_n5669 = n2183 & new_n5667;
  assign new_n5670 = n2182 & new_n5667;
  assign new_n5671 = n2181 & new_n5667;
  assign new_n5672 = n2180 & new_n5667;
  assign new_n5673 = n2179 & new_n5667;
  assign new_n5674 = n2178 & new_n5667;
  assign new_n5675 = n2177 & new_n5667;
  assign new_n5676 = new_n5427 & new_n5484;
  assign new_n5677 = new_n5434 & new_n5676;
  assign new_n5678 = new_n5430 & new_n5676;
  assign new_n5679 = ~new_n5677 & ~new_n5678;
  assign new_n5680 = new_n5438 & new_n5676;
  assign new_n5681 = ~new_n5680 & new_n5679;
  assign new_n5682 = n2240 & new_n5681;
  assign new_n5683 = n2239 & new_n5681;
  assign new_n5684 = n2238 & new_n5681;
  assign new_n5685 = n2237 & new_n5681;
  assign new_n5686 = n2236 & new_n5681;
  assign new_n5687 = n2235 & new_n5681;
  assign new_n5688 = n2234 & new_n5681;
  assign new_n5689 = n2233 & new_n5681;
  assign new_n5690 = new_n5500 & new_n5676;
  assign new_n5691 = ~new_n5690 & new_n5679;
  assign new_n5692 = n2232 & new_n5691;
  assign new_n5693 = n2231 & new_n5691;
  assign new_n5694 = n2230 & new_n5691;
  assign new_n5695 = n2229 & new_n5691;
  assign new_n5696 = n2228 & new_n5691;
  assign new_n5697 = n2227 & new_n5691;
  assign new_n5698 = n2226 & new_n5691;
  assign new_n5699 = n2225 & new_n5691;
  assign new_n5700 = new_n5433 & new_n5676;
  assign new_n5701 = ~new_n5678 & ~new_n5700;
  assign new_n5702 = new_n5513 & new_n5676;
  assign new_n5703 = ~new_n5702 & new_n5701;
  assign new_n5704 = n2224 & new_n5703;
  assign new_n5705 = n2223 & new_n5703;
  assign new_n5706 = n2222 & new_n5703;
  assign new_n5707 = n2221 & new_n5703;
  assign new_n5708 = n2220 & new_n5703;
  assign new_n5709 = n2219 & new_n5703;
  assign new_n5710 = n2218 & new_n5703;
  assign new_n5711 = n2217 & new_n5703;
  assign new_n5712 = new_n5524 & new_n5676;
  assign new_n5713 = ~new_n5712 & new_n5701;
  assign new_n5714 = n2216 & new_n5713;
  assign new_n5715 = n2215 & new_n5713;
  assign new_n5716 = n2214 & new_n5713;
  assign new_n5717 = n2213 & new_n5713;
  assign new_n5718 = n2212 & new_n5713;
  assign new_n5719 = n2211 & new_n5713;
  assign new_n5720 = n2210 & new_n5713;
  assign new_n5721 = n2209 & new_n5713;
  assign new_n5722 = new_n5427 & new_n5536;
  assign new_n5723 = new_n5434 & new_n5722;
  assign new_n5724 = new_n5430 & new_n5722;
  assign new_n5725 = ~new_n5723 & ~new_n5724;
  assign new_n5726 = new_n5438 & new_n5722;
  assign new_n5727 = ~new_n5726 & new_n5725;
  assign new_n5728 = n2272 & new_n5727;
  assign new_n5729 = n2271 & new_n5727;
  assign new_n5730 = n2270 & new_n5727;
  assign new_n5731 = n2269 & new_n5727;
  assign new_n5732 = n2268 & new_n5727;
  assign new_n5733 = n2267 & new_n5727;
  assign new_n5734 = n2266 & new_n5727;
  assign new_n5735 = n2265 & new_n5727;
  assign new_n5736 = new_n5500 & new_n5722;
  assign new_n5737 = ~new_n5736 & new_n5725;
  assign new_n5738 = n2264 & new_n5737;
  assign new_n5739 = n2263 & new_n5737;
  assign new_n5740 = n2262 & new_n5737;
  assign new_n5741 = n2261 & new_n5737;
  assign new_n5742 = n2260 & new_n5737;
  assign new_n5743 = n2259 & new_n5737;
  assign new_n5744 = n2258 & new_n5737;
  assign new_n5745 = n2257 & new_n5737;
  assign new_n5746 = new_n5433 & new_n5722;
  assign new_n5747 = ~new_n5724 & ~new_n5746;
  assign new_n5748 = new_n5513 & new_n5722;
  assign new_n5749 = ~new_n5748 & new_n5747;
  assign new_n5750 = n2256 & new_n5749;
  assign new_n5751 = n2255 & new_n5749;
  assign new_n5752 = n2254 & new_n5749;
  assign new_n5753 = n2253 & new_n5749;
  assign new_n5754 = n2252 & new_n5749;
  assign new_n5755 = n2251 & new_n5749;
  assign new_n5756 = n2250 & new_n5749;
  assign new_n5757 = n2249 & new_n5749;
  assign new_n5758 = new_n5524 & new_n5722;
  assign new_n5759 = ~new_n5758 & new_n5747;
  assign new_n5760 = n2248 & new_n5759;
  assign new_n5761 = n2247 & new_n5759;
  assign new_n5762 = n2246 & new_n5759;
  assign new_n5763 = n2245 & new_n5759;
  assign new_n5764 = n2244 & new_n5759;
  assign new_n5765 = n2243 & new_n5759;
  assign new_n5766 = n2242 & new_n5759;
  assign new_n5767 = n2241 & new_n5759;
  assign new_n5768 = new_n5246 & new_n5427;
  assign new_n5769 = new_n5434 & new_n5768;
  assign new_n5770 = new_n5430 & new_n5768;
  assign new_n5771 = ~new_n5769 & ~new_n5770;
  assign new_n5772 = new_n5438 & new_n5768;
  assign new_n5773 = ~new_n5772 & new_n5771;
  assign new_n5774 = n2304 & new_n5773;
  assign new_n5775 = n2303 & new_n5773;
  assign new_n5776 = n2302 & new_n5773;
  assign new_n5777 = n2301 & new_n5773;
  assign new_n5778 = n2300 & new_n5773;
  assign new_n5779 = n2299 & new_n5773;
  assign new_n5780 = n2298 & new_n5773;
  assign new_n5781 = n2297 & new_n5773;
  assign new_n5782 = new_n5500 & new_n5768;
  assign new_n5783 = ~new_n5782 & new_n5771;
  assign new_n5784 = n2296 & new_n5783;
  assign new_n5785 = n2295 & new_n5783;
  assign new_n5786 = n2294 & new_n5783;
  assign new_n5787 = n2293 & new_n5783;
  assign new_n5788 = n2292 & new_n5783;
  assign new_n5789 = n2291 & new_n5783;
  assign new_n5790 = n2290 & new_n5783;
  assign new_n5791 = n2289 & new_n5783;
  assign new_n5792 = new_n5433 & new_n5768;
  assign new_n5793 = ~new_n5770 & ~new_n5792;
  assign new_n5794 = new_n5513 & new_n5768;
  assign new_n5795 = ~new_n5794 & new_n5793;
  assign new_n5796 = n2288 & new_n5795;
  assign new_n5797 = n2287 & new_n5795;
  assign new_n5798 = n2286 & new_n5795;
  assign new_n5799 = n2285 & new_n5795;
  assign new_n5800 = n2284 & new_n5795;
  assign new_n5801 = n2283 & new_n5795;
  assign new_n5802 = n2282 & new_n5795;
  assign new_n5803 = n2281 & new_n5795;
  assign new_n5804 = new_n5524 & new_n5768;
  assign new_n5805 = ~new_n5804 & new_n5793;
  assign new_n5806 = n2280 & new_n5805;
  assign new_n5807 = n2279 & new_n5805;
  assign new_n5808 = n2278 & new_n5805;
  assign new_n5809 = n2277 & new_n5805;
  assign new_n5810 = n2276 & new_n5805;
  assign new_n5811 = n2275 & new_n5805;
  assign new_n5812 = n2274 & new_n5805;
  assign new_n5813 = n2273 & new_n5805;
  assign new_n5814 = ~new_n5011 & new_n5139;
  assign new_n5815 = new_n5031 & new_n5814;
  assign new_n5816 = new_n5815 ^ new_n5814;
  assign new_n5817 = new_n5424 & new_n5816;
  assign new_n5818 = new_n5434 & new_n5817;
  assign new_n5819 = new_n5430 & new_n5817;
  assign new_n5820 = ~new_n5818 & ~new_n5819;
  assign new_n5821 = new_n5438 & new_n5817;
  assign new_n5822 = ~new_n5821 & new_n5820;
  assign new_n5823 = n2336 & new_n5822;
  assign new_n5824 = n2335 & new_n5822;
  assign new_n5825 = n2334 & new_n5822;
  assign new_n5826 = n2333 & new_n5822;
  assign new_n5827 = n2332 & new_n5822;
  assign new_n5828 = n2331 & new_n5822;
  assign new_n5829 = n2330 & new_n5822;
  assign new_n5830 = n2329 & new_n5822;
  assign new_n5831 = new_n5500 & new_n5817;
  assign new_n5832 = ~new_n5831 & new_n5820;
  assign new_n5833 = n2328 & new_n5832;
  assign new_n5834 = n2327 & new_n5832;
  assign new_n5835 = n2326 & new_n5832;
  assign new_n5836 = n2325 & new_n5832;
  assign new_n5837 = n2324 & new_n5832;
  assign new_n5838 = n2323 & new_n5832;
  assign new_n5839 = n2322 & new_n5832;
  assign new_n5840 = n2321 & new_n5832;
  assign new_n5841 = new_n5433 & new_n5817;
  assign new_n5842 = ~new_n5819 & ~new_n5841;
  assign new_n5843 = new_n5513 & new_n5817;
  assign new_n5844 = ~new_n5843 & new_n5842;
  assign new_n5845 = n2320 & new_n5844;
  assign new_n5846 = n2319 & new_n5844;
  assign new_n5847 = n2318 & new_n5844;
  assign new_n5848 = n2317 & new_n5844;
  assign new_n5849 = n2316 & new_n5844;
  assign new_n5850 = n2315 & new_n5844;
  assign new_n5851 = n2314 & new_n5844;
  assign new_n5852 = n2313 & new_n5844;
  assign new_n5853 = new_n5524 & new_n5817;
  assign new_n5854 = ~new_n5853 & new_n5842;
  assign new_n5855 = n2312 & new_n5854;
  assign new_n5856 = n2311 & new_n5854;
  assign new_n5857 = n2310 & new_n5854;
  assign new_n5858 = n2309 & new_n5854;
  assign new_n5859 = n2308 & new_n5854;
  assign new_n5860 = n2307 & new_n5854;
  assign new_n5861 = n2306 & new_n5854;
  assign new_n5862 = n2305 & new_n5854;
  assign new_n5863 = new_n5485 & new_n5816;
  assign new_n5864 = new_n5434 & new_n5863;
  assign new_n5865 = new_n5430 & new_n5863;
  assign new_n5866 = ~new_n5864 & ~new_n5865;
  assign new_n5867 = new_n5438 & new_n5863;
  assign new_n5868 = ~new_n5867 & new_n5866;
  assign new_n5869 = n2368 & new_n5868;
  assign new_n5870 = n2367 & new_n5868;
  assign new_n5871 = n2366 & new_n5868;
  assign new_n5872 = n2365 & new_n5868;
  assign new_n5873 = n2364 & new_n5868;
  assign new_n5874 = n2363 & new_n5868;
  assign new_n5875 = n2362 & new_n5868;
  assign new_n5876 = n2361 & new_n5868;
  assign new_n5877 = new_n5500 & new_n5863;
  assign new_n5878 = ~new_n5877 & new_n5866;
  assign new_n5879 = n2360 & new_n5878;
  assign new_n5880 = n2359 & new_n5878;
  assign new_n5881 = n2358 & new_n5878;
  assign new_n5882 = n2357 & new_n5878;
  assign new_n5883 = n2356 & new_n5878;
  assign new_n5884 = n2355 & new_n5878;
  assign new_n5885 = n2354 & new_n5878;
  assign new_n5886 = n2353 & new_n5878;
  assign new_n5887 = new_n5433 & new_n5863;
  assign new_n5888 = ~new_n5865 & ~new_n5887;
  assign new_n5889 = new_n5513 & new_n5863;
  assign new_n5890 = ~new_n5889 & new_n5888;
  assign new_n5891 = n2352 & new_n5890;
  assign new_n5892 = n2351 & new_n5890;
  assign new_n5893 = n2350 & new_n5890;
  assign new_n5894 = n2349 & new_n5890;
  assign new_n5895 = n2348 & new_n5890;
  assign new_n5896 = n2347 & new_n5890;
  assign new_n5897 = n2346 & new_n5890;
  assign new_n5898 = n2345 & new_n5890;
  assign new_n5899 = new_n5524 & new_n5863;
  assign new_n5900 = ~new_n5899 & new_n5888;
  assign new_n5901 = n2344 & new_n5900;
  assign new_n5902 = n2343 & new_n5900;
  assign new_n5903 = n2342 & new_n5900;
  assign new_n5904 = n2341 & new_n5900;
  assign new_n5905 = n2340 & new_n5900;
  assign new_n5906 = n2339 & new_n5900;
  assign new_n5907 = n2338 & new_n5900;
  assign new_n5908 = n2337 & new_n5900;
  assign new_n5909 = new_n5537 & new_n5816;
  assign new_n5910 = new_n5434 & new_n5909;
  assign new_n5911 = new_n5430 & new_n5909;
  assign new_n5912 = ~new_n5910 & ~new_n5911;
  assign new_n5913 = new_n5438 & new_n5909;
  assign new_n5914 = ~new_n5913 & new_n5912;
  assign new_n5915 = n2400 & new_n5914;
  assign new_n5916 = n2399 & new_n5914;
  assign new_n5917 = n2398 & new_n5914;
  assign new_n5918 = n2397 & new_n5914;
  assign new_n5919 = n2396 & new_n5914;
  assign new_n5920 = n2395 & new_n5914;
  assign new_n5921 = n2394 & new_n5914;
  assign new_n5922 = n2393 & new_n5914;
  assign new_n5923 = new_n5500 & new_n5909;
  assign new_n5924 = ~new_n5923 & new_n5912;
  assign new_n5925 = n2392 & new_n5924;
  assign new_n5926 = n2391 & new_n5924;
  assign new_n5927 = n2390 & new_n5924;
  assign new_n5928 = n2389 & new_n5924;
  assign new_n5929 = n2388 & new_n5924;
  assign new_n5930 = n2387 & new_n5924;
  assign new_n5931 = n2386 & new_n5924;
  assign new_n5932 = n2385 & new_n5924;
  assign new_n5933 = new_n5433 & new_n5909;
  assign new_n5934 = ~new_n5911 & ~new_n5933;
  assign new_n5935 = new_n5513 & new_n5909;
  assign new_n5936 = ~new_n5935 & new_n5934;
  assign new_n5937 = n2384 & new_n5936;
  assign new_n5938 = n2383 & new_n5936;
  assign new_n5939 = n2382 & new_n5936;
  assign new_n5940 = n2381 & new_n5936;
  assign new_n5941 = n2380 & new_n5936;
  assign new_n5942 = n2379 & new_n5936;
  assign new_n5943 = n2378 & new_n5936;
  assign new_n5944 = n2377 & new_n5936;
  assign new_n5945 = new_n5524 & new_n5909;
  assign new_n5946 = ~new_n5945 & new_n5934;
  assign new_n5947 = n2376 & new_n5946;
  assign new_n5948 = n2375 & new_n5946;
  assign new_n5949 = n2374 & new_n5946;
  assign new_n5950 = n2373 & new_n5946;
  assign new_n5951 = n2372 & new_n5946;
  assign new_n5952 = n2371 & new_n5946;
  assign new_n5953 = n2370 & new_n5946;
  assign new_n5954 = n2369 & new_n5946;
  assign new_n5955 = new_n5245 & new_n5816;
  assign new_n5956 = new_n5434 & new_n5955;
  assign new_n5957 = new_n5430 & new_n5955;
  assign new_n5958 = ~new_n5956 & ~new_n5957;
  assign new_n5959 = new_n5438 & new_n5955;
  assign new_n5960 = ~new_n5959 & new_n5958;
  assign new_n5961 = n2432 & new_n5960;
  assign new_n5962 = n2431 & new_n5960;
  assign new_n5963 = n2430 & new_n5960;
  assign new_n5964 = n2429 & new_n5960;
  assign new_n5965 = n2428 & new_n5960;
  assign new_n5966 = n2427 & new_n5960;
  assign new_n5967 = n2426 & new_n5960;
  assign new_n5968 = n2425 & new_n5960;
  assign new_n5969 = new_n5500 & new_n5955;
  assign new_n5970 = ~new_n5969 & new_n5958;
  assign new_n5971 = n2424 & new_n5970;
  assign new_n5972 = n2423 & new_n5970;
  assign new_n5973 = n2422 & new_n5970;
  assign new_n5974 = n2421 & new_n5970;
  assign new_n5975 = n2420 & new_n5970;
  assign new_n5976 = n2419 & new_n5970;
  assign new_n5977 = n2418 & new_n5970;
  assign new_n5978 = n2417 & new_n5970;
  assign new_n5979 = new_n5433 & new_n5955;
  assign new_n5980 = ~new_n5957 & ~new_n5979;
  assign new_n5981 = new_n5513 & new_n5955;
  assign new_n5982 = ~new_n5981 & new_n5980;
  assign new_n5983 = n2416 & new_n5982;
  assign new_n5984 = n2415 & new_n5982;
  assign new_n5985 = n2414 & new_n5982;
  assign new_n5986 = n2413 & new_n5982;
  assign new_n5987 = n2412 & new_n5982;
  assign new_n5988 = n2411 & new_n5982;
  assign new_n5989 = n2410 & new_n5982;
  assign new_n5990 = n2409 & new_n5982;
  assign new_n5991 = new_n5524 & new_n5955;
  assign new_n5992 = ~new_n5991 & new_n5980;
  assign new_n5993 = n2408 & new_n5992;
  assign new_n5994 = n2407 & new_n5992;
  assign new_n5995 = n2406 & new_n5992;
  assign new_n5996 = n2405 & new_n5992;
  assign new_n5997 = n2404 & new_n5992;
  assign new_n5998 = n2403 & new_n5992;
  assign new_n5999 = n2402 & new_n5992;
  assign new_n6000 = n2401 & new_n5992;
  assign new_n6001 = new_n5423 & new_n5816;
  assign new_n6002 = new_n5434 & new_n6001;
  assign new_n6003 = new_n5430 & new_n6001;
  assign new_n6004 = ~new_n6002 & ~new_n6003;
  assign new_n6005 = new_n5438 & new_n6001;
  assign new_n6006 = ~new_n6005 & new_n6004;
  assign new_n6007 = n2464 & new_n6006;
  assign new_n6008 = n2463 & new_n6006;
  assign new_n6009 = n2462 & new_n6006;
  assign new_n6010 = n2461 & new_n6006;
  assign new_n6011 = n2460 & new_n6006;
  assign new_n6012 = n2459 & new_n6006;
  assign new_n6013 = n2458 & new_n6006;
  assign new_n6014 = n2457 & new_n6006;
  assign new_n6015 = new_n5500 & new_n6001;
  assign new_n6016 = ~new_n6015 & new_n6004;
  assign new_n6017 = n2456 & new_n6016;
  assign new_n6018 = n2455 & new_n6016;
  assign new_n6019 = n2454 & new_n6016;
  assign new_n6020 = n2453 & new_n6016;
  assign new_n6021 = n2452 & new_n6016;
  assign new_n6022 = n2451 & new_n6016;
  assign new_n6023 = n2450 & new_n6016;
  assign new_n6024 = n2449 & new_n6016;
  assign new_n6025 = new_n5433 & new_n6001;
  assign new_n6026 = ~new_n6003 & ~new_n6025;
  assign new_n6027 = new_n5513 & new_n6001;
  assign new_n6028 = ~new_n6027 & new_n6026;
  assign new_n6029 = n2448 & new_n6028;
  assign new_n6030 = n2447 & new_n6028;
  assign new_n6031 = n2446 & new_n6028;
  assign new_n6032 = n2445 & new_n6028;
  assign new_n6033 = n2444 & new_n6028;
  assign new_n6034 = n2443 & new_n6028;
  assign new_n6035 = n2442 & new_n6028;
  assign new_n6036 = n2441 & new_n6028;
  assign new_n6037 = new_n5524 & new_n6001;
  assign new_n6038 = ~new_n6037 & new_n6026;
  assign new_n6039 = n2440 & new_n6038;
  assign new_n6040 = n2439 & new_n6038;
  assign new_n6041 = n2438 & new_n6038;
  assign new_n6042 = n2437 & new_n6038;
  assign new_n6043 = n2436 & new_n6038;
  assign new_n6044 = n2435 & new_n6038;
  assign new_n6045 = n2434 & new_n6038;
  assign new_n6046 = n2433 & new_n6038;
  assign new_n6047 = new_n5484 & new_n5816;
  assign new_n6048 = new_n5434 & new_n6047;
  assign new_n6049 = new_n5430 & new_n6047;
  assign new_n6050 = ~new_n6048 & ~new_n6049;
  assign new_n6051 = new_n5438 & new_n6047;
  assign new_n6052 = ~new_n6051 & new_n6050;
  assign new_n6053 = n2496 & new_n6052;
  assign new_n6054 = n2495 & new_n6052;
  assign new_n6055 = n2494 & new_n6052;
  assign new_n6056 = n2493 & new_n6052;
  assign new_n6057 = n2492 & new_n6052;
  assign new_n6058 = n2491 & new_n6052;
  assign new_n6059 = n2490 & new_n6052;
  assign new_n6060 = n2489 & new_n6052;
  assign new_n6061 = new_n5500 & new_n6047;
  assign new_n6062 = ~new_n6061 & new_n6050;
  assign new_n6063 = n2488 & new_n6062;
  assign new_n6064 = n2487 & new_n6062;
  assign new_n6065 = n2486 & new_n6062;
  assign new_n6066 = n2485 & new_n6062;
  assign new_n6067 = n2484 & new_n6062;
  assign new_n6068 = n2483 & new_n6062;
  assign new_n6069 = n2482 & new_n6062;
  assign new_n6070 = n2481 & new_n6062;
  assign new_n6071 = new_n5433 & new_n6047;
  assign new_n6072 = ~new_n6049 & ~new_n6071;
  assign new_n6073 = new_n5513 & new_n6047;
  assign new_n6074 = ~new_n6073 & new_n6072;
  assign new_n6075 = n2480 & new_n6074;
  assign new_n6076 = n2479 & new_n6074;
  assign new_n6077 = n2478 & new_n6074;
  assign new_n6078 = n2477 & new_n6074;
  assign new_n6079 = n2476 & new_n6074;
  assign new_n6080 = n2475 & new_n6074;
  assign new_n6081 = n2474 & new_n6074;
  assign new_n6082 = n2473 & new_n6074;
  assign new_n6083 = new_n5524 & new_n6047;
  assign new_n6084 = ~new_n6083 & new_n6072;
  assign new_n6085 = n2472 & new_n6084;
  assign new_n6086 = n2471 & new_n6084;
  assign new_n6087 = n2470 & new_n6084;
  assign new_n6088 = n2469 & new_n6084;
  assign new_n6089 = n2468 & new_n6084;
  assign new_n6090 = n2467 & new_n6084;
  assign new_n6091 = n2466 & new_n6084;
  assign new_n6092 = n2465 & new_n6084;
  assign new_n6093 = new_n5536 & new_n5816;
  assign new_n6094 = new_n5434 & new_n6093;
  assign new_n6095 = new_n5430 & new_n6093;
  assign new_n6096 = ~new_n6094 & ~new_n6095;
  assign new_n6097 = new_n5438 & new_n6093;
  assign new_n6098 = ~new_n6097 & new_n6096;
  assign new_n6099 = n2528 & new_n6098;
  assign new_n6100 = n2527 & new_n6098;
  assign new_n6101 = n2526 & new_n6098;
  assign new_n6102 = n2525 & new_n6098;
  assign new_n6103 = n2524 & new_n6098;
  assign new_n6104 = n2523 & new_n6098;
  assign new_n6105 = n2522 & new_n6098;
  assign new_n6106 = n2521 & new_n6098;
  assign new_n6107 = new_n5500 & new_n6093;
  assign new_n6108 = ~new_n6107 & new_n6096;
  assign new_n6109 = n2520 & new_n6108;
  assign new_n6110 = n2519 & new_n6108;
  assign new_n6111 = n2518 & new_n6108;
  assign new_n6112 = n2517 & new_n6108;
  assign new_n6113 = n2516 & new_n6108;
  assign new_n6114 = n2515 & new_n6108;
  assign new_n6115 = n2514 & new_n6108;
  assign new_n6116 = n2513 & new_n6108;
  assign new_n6117 = new_n5433 & new_n6093;
  assign new_n6118 = ~new_n6095 & ~new_n6117;
  assign new_n6119 = new_n5513 & new_n6093;
  assign new_n6120 = ~new_n6119 & new_n6118;
  assign new_n6121 = n2512 & new_n6120;
  assign new_n6122 = n2511 & new_n6120;
  assign new_n6123 = n2510 & new_n6120;
  assign new_n6124 = n2509 & new_n6120;
  assign new_n6125 = n2508 & new_n6120;
  assign new_n6126 = n2507 & new_n6120;
  assign new_n6127 = n2506 & new_n6120;
  assign new_n6128 = n2505 & new_n6120;
  assign new_n6129 = new_n5524 & new_n6093;
  assign new_n6130 = ~new_n6129 & new_n6118;
  assign new_n6131 = n2504 & new_n6130;
  assign new_n6132 = n2503 & new_n6130;
  assign new_n6133 = n2502 & new_n6130;
  assign new_n6134 = n2501 & new_n6130;
  assign new_n6135 = n2500 & new_n6130;
  assign new_n6136 = n2499 & new_n6130;
  assign new_n6137 = n2498 & new_n6130;
  assign new_n6138 = n2497 & new_n6130;
  assign new_n6139 = new_n5246 & new_n5816;
  assign new_n6140 = new_n5434 & new_n6139;
  assign new_n6141 = new_n5430 & new_n6139;
  assign new_n6142 = ~new_n6140 & ~new_n6141;
  assign new_n6143 = new_n5438 & new_n6139;
  assign new_n6144 = ~new_n6143 & new_n6142;
  assign new_n6145 = n2560 & new_n6144;
  assign new_n6146 = n2559 & new_n6144;
  assign new_n6147 = n2558 & new_n6144;
  assign new_n6148 = n2557 & new_n6144;
  assign new_n6149 = n2556 & new_n6144;
  assign new_n6150 = n2555 & new_n6144;
  assign new_n6151 = n2554 & new_n6144;
  assign new_n6152 = n2553 & new_n6144;
  assign new_n6153 = new_n5500 & new_n6139;
  assign new_n6154 = ~new_n6153 & new_n6142;
  assign new_n6155 = n2552 & new_n6154;
  assign new_n6156 = n2551 & new_n6154;
  assign new_n6157 = n2550 & new_n6154;
  assign new_n6158 = n2549 & new_n6154;
  assign new_n6159 = n2548 & new_n6154;
  assign new_n6160 = n2547 & new_n6154;
  assign new_n6161 = n2546 & new_n6154;
  assign new_n6162 = n2545 & new_n6154;
  assign new_n6163 = new_n5433 & new_n6139;
  assign new_n6164 = ~new_n6141 & ~new_n6163;
  assign new_n6165 = new_n5513 & new_n6139;
  assign new_n6166 = ~new_n6165 & new_n6164;
  assign new_n6167 = n2544 & new_n6166;
  assign new_n6168 = n2543 & new_n6166;
  assign new_n6169 = n2542 & new_n6166;
  assign new_n6170 = n2541 & new_n6166;
  assign new_n6171 = n2540 & new_n6166;
  assign new_n6172 = n2539 & new_n6166;
  assign new_n6173 = n2538 & new_n6166;
  assign new_n6174 = n2537 & new_n6166;
  assign new_n6175 = new_n5524 & new_n6139;
  assign new_n6176 = ~new_n6175 & new_n6164;
  assign new_n6177 = n2536 & new_n6176;
  assign new_n6178 = n2535 & new_n6176;
  assign new_n6179 = n2534 & new_n6176;
  assign new_n6180 = n2533 & new_n6176;
  assign new_n6181 = n2532 & new_n6176;
  assign new_n6182 = n2531 & new_n6176;
  assign new_n6183 = n2530 & new_n6176;
  assign new_n6184 = n2529 & new_n6176;
  assign new_n6185 = ~new_n5139 & new_n5011;
  assign new_n6186 = new_n5031 & new_n6185;
  assign new_n6187 = new_n6186 ^ new_n6185;
  assign new_n6188 = new_n5424 & new_n6187;
  assign new_n6189 = new_n5434 & new_n6188;
  assign new_n6190 = new_n5430 & new_n6188;
  assign new_n6191 = ~new_n6189 & ~new_n6190;
  assign new_n6192 = new_n5438 & new_n6188;
  assign new_n6193 = ~new_n6192 & new_n6191;
  assign new_n6194 = n2592 & new_n6193;
  assign new_n6195 = n2591 & new_n6193;
  assign new_n6196 = n2590 & new_n6193;
  assign new_n6197 = n2589 & new_n6193;
  assign new_n6198 = n2588 & new_n6193;
  assign new_n6199 = n2587 & new_n6193;
  assign new_n6200 = n2586 & new_n6193;
  assign new_n6201 = n2585 & new_n6193;
  assign new_n6202 = new_n5500 & new_n6188;
  assign new_n6203 = ~new_n6202 & new_n6191;
  assign new_n6204 = n2584 & new_n6203;
  assign new_n6205 = n2583 & new_n6203;
  assign new_n6206 = n2582 & new_n6203;
  assign new_n6207 = n2581 & new_n6203;
  assign new_n6208 = n2580 & new_n6203;
  assign new_n6209 = n2579 & new_n6203;
  assign new_n6210 = n2578 & new_n6203;
  assign new_n6211 = n2577 & new_n6203;
  assign new_n6212 = new_n5433 & new_n6188;
  assign new_n6213 = ~new_n6190 & ~new_n6212;
  assign new_n6214 = new_n5513 & new_n6188;
  assign new_n6215 = ~new_n6214 & new_n6213;
  assign new_n6216 = n2576 & new_n6215;
  assign new_n6217 = n2575 & new_n6215;
  assign new_n6218 = n2574 & new_n6215;
  assign new_n6219 = n2573 & new_n6215;
  assign new_n6220 = n2572 & new_n6215;
  assign new_n6221 = n2571 & new_n6215;
  assign new_n6222 = n2570 & new_n6215;
  assign new_n6223 = n2569 & new_n6215;
  assign new_n6224 = new_n5524 & new_n6188;
  assign new_n6225 = ~new_n6224 & new_n6213;
  assign new_n6226 = n2568 & new_n6225;
  assign new_n6227 = n2567 & new_n6225;
  assign new_n6228 = n2566 & new_n6225;
  assign new_n6229 = n2565 & new_n6225;
  assign new_n6230 = n2564 & new_n6225;
  assign new_n6231 = n2563 & new_n6225;
  assign new_n6232 = n2562 & new_n6225;
  assign new_n6233 = n2561 & new_n6225;
  assign new_n6234 = new_n5485 & new_n6187;
  assign new_n6235 = new_n5434 & new_n6234;
  assign new_n6236 = new_n5430 & new_n6234;
  assign new_n6237 = ~new_n6235 & ~new_n6236;
  assign new_n6238 = new_n5438 & new_n6234;
  assign new_n6239 = ~new_n6238 & new_n6237;
  assign new_n6240 = n2624 & new_n6239;
  assign new_n6241 = n2623 & new_n6239;
  assign new_n6242 = n2622 & new_n6239;
  assign new_n6243 = n2621 & new_n6239;
  assign new_n6244 = n2620 & new_n6239;
  assign new_n6245 = n2619 & new_n6239;
  assign new_n6246 = n2618 & new_n6239;
  assign new_n6247 = n2617 & new_n6239;
  assign new_n6248 = new_n5500 & new_n6234;
  assign new_n6249 = ~new_n6248 & new_n6237;
  assign new_n6250 = n2616 & new_n6249;
  assign new_n6251 = n2615 & new_n6249;
  assign new_n6252 = n2614 & new_n6249;
  assign new_n6253 = n2613 & new_n6249;
  assign new_n6254 = n2612 & new_n6249;
  assign new_n6255 = n2611 & new_n6249;
  assign new_n6256 = n2610 & new_n6249;
  assign new_n6257 = n2609 & new_n6249;
  assign new_n6258 = new_n5433 & new_n6234;
  assign new_n6259 = ~new_n6236 & ~new_n6258;
  assign new_n6260 = new_n5513 & new_n6234;
  assign new_n6261 = ~new_n6260 & new_n6259;
  assign new_n6262 = n2608 & new_n6261;
  assign new_n6263 = n2607 & new_n6261;
  assign new_n6264 = n2606 & new_n6261;
  assign new_n6265 = n2605 & new_n6261;
  assign new_n6266 = n2604 & new_n6261;
  assign new_n6267 = n2603 & new_n6261;
  assign new_n6268 = n2602 & new_n6261;
  assign new_n6269 = n2601 & new_n6261;
  assign new_n6270 = new_n5524 & new_n6234;
  assign new_n6271 = ~new_n6270 & new_n6259;
  assign new_n6272 = n2600 & new_n6271;
  assign new_n6273 = n2599 & new_n6271;
  assign new_n6274 = n2598 & new_n6271;
  assign new_n6275 = n2597 & new_n6271;
  assign new_n6276 = n2596 & new_n6271;
  assign new_n6277 = n2595 & new_n6271;
  assign new_n6278 = n2594 & new_n6271;
  assign new_n6279 = n2593 & new_n6271;
  assign new_n6280 = new_n5537 & new_n6187;
  assign new_n6281 = new_n5434 & new_n6280;
  assign new_n6282 = new_n5430 & new_n6280;
  assign new_n6283 = ~new_n6281 & ~new_n6282;
  assign new_n6284 = new_n5438 & new_n6280;
  assign new_n6285 = ~new_n6284 & new_n6283;
  assign new_n6286 = n2656 & new_n6285;
  assign new_n6287 = n2655 & new_n6285;
  assign new_n6288 = n2654 & new_n6285;
  assign new_n6289 = n2653 & new_n6285;
  assign new_n6290 = n2652 & new_n6285;
  assign new_n6291 = n2651 & new_n6285;
  assign new_n6292 = n2650 & new_n6285;
  assign new_n6293 = n2649 & new_n6285;
  assign new_n6294 = new_n5500 & new_n6280;
  assign new_n6295 = ~new_n6294 & new_n6283;
  assign new_n6296 = n2648 & new_n6295;
  assign new_n6297 = n2647 & new_n6295;
  assign new_n6298 = n2646 & new_n6295;
  assign new_n6299 = n2645 & new_n6295;
  assign new_n6300 = n2644 & new_n6295;
  assign new_n6301 = n2643 & new_n6295;
  assign new_n6302 = n2642 & new_n6295;
  assign new_n6303 = n2641 & new_n6295;
  assign new_n6304 = new_n5433 & new_n6280;
  assign new_n6305 = ~new_n6282 & ~new_n6304;
  assign new_n6306 = new_n5513 & new_n6280;
  assign new_n6307 = ~new_n6306 & new_n6305;
  assign new_n6308 = n2640 & new_n6307;
  assign new_n6309 = n2639 & new_n6307;
  assign new_n6310 = n2638 & new_n6307;
  assign new_n6311 = n2637 & new_n6307;
  assign new_n6312 = n2636 & new_n6307;
  assign new_n6313 = n2635 & new_n6307;
  assign new_n6314 = n2634 & new_n6307;
  assign new_n6315 = n2633 & new_n6307;
  assign new_n6316 = new_n5524 & new_n6280;
  assign new_n6317 = ~new_n6316 & new_n6305;
  assign new_n6318 = n2632 & new_n6317;
  assign new_n6319 = n2631 & new_n6317;
  assign new_n6320 = n2630 & new_n6317;
  assign new_n6321 = n2629 & new_n6317;
  assign new_n6322 = n2628 & new_n6317;
  assign new_n6323 = n2627 & new_n6317;
  assign new_n6324 = n2626 & new_n6317;
  assign new_n6325 = n2625 & new_n6317;
  assign new_n6326 = new_n5245 & new_n6187;
  assign new_n6327 = new_n5434 & new_n6326;
  assign new_n6328 = new_n5430 & new_n6326;
  assign new_n6329 = ~new_n6327 & ~new_n6328;
  assign new_n6330 = new_n5438 & new_n6326;
  assign new_n6331 = ~new_n6330 & new_n6329;
  assign new_n6332 = n2688 & new_n6331;
  assign new_n6333 = n2687 & new_n6331;
  assign new_n6334 = n2686 & new_n6331;
  assign new_n6335 = n2685 & new_n6331;
  assign new_n6336 = n2684 & new_n6331;
  assign new_n6337 = n2683 & new_n6331;
  assign new_n6338 = n2682 & new_n6331;
  assign new_n6339 = n2681 & new_n6331;
  assign new_n6340 = new_n5500 & new_n6326;
  assign new_n6341 = ~new_n6340 & new_n6329;
  assign new_n6342 = n2680 & new_n6341;
  assign new_n6343 = n2679 & new_n6341;
  assign new_n6344 = n2678 & new_n6341;
  assign new_n6345 = n2677 & new_n6341;
  assign new_n6346 = n2676 & new_n6341;
  assign new_n6347 = n2675 & new_n6341;
  assign new_n6348 = n2674 & new_n6341;
  assign new_n6349 = n2673 & new_n6341;
  assign new_n6350 = new_n5433 & new_n6326;
  assign new_n6351 = ~new_n6328 & ~new_n6350;
  assign new_n6352 = new_n5513 & new_n6326;
  assign new_n6353 = ~new_n6352 & new_n6351;
  assign new_n6354 = n2672 & new_n6353;
  assign new_n6355 = n2671 & new_n6353;
  assign new_n6356 = n2670 & new_n6353;
  assign new_n6357 = n2669 & new_n6353;
  assign new_n6358 = n2668 & new_n6353;
  assign new_n6359 = n2667 & new_n6353;
  assign new_n6360 = n2666 & new_n6353;
  assign new_n6361 = n2665 & new_n6353;
  assign new_n6362 = new_n5524 & new_n6326;
  assign new_n6363 = ~new_n6362 & new_n6351;
  assign new_n6364 = n2664 & new_n6363;
  assign new_n6365 = n2663 & new_n6363;
  assign new_n6366 = n2662 & new_n6363;
  assign new_n6367 = n2661 & new_n6363;
  assign new_n6368 = n2660 & new_n6363;
  assign new_n6369 = n2659 & new_n6363;
  assign new_n6370 = n2658 & new_n6363;
  assign new_n6371 = n2657 & new_n6363;
  assign new_n6372 = new_n5423 & new_n6187;
  assign new_n6373 = new_n5434 & new_n6372;
  assign new_n6374 = new_n5430 & new_n6372;
  assign new_n6375 = ~new_n6373 & ~new_n6374;
  assign new_n6376 = new_n5438 & new_n6372;
  assign new_n6377 = ~new_n6376 & new_n6375;
  assign new_n6378 = n2720 & new_n6377;
  assign new_n6379 = n2719 & new_n6377;
  assign new_n6380 = n2718 & new_n6377;
  assign new_n6381 = n2717 & new_n6377;
  assign new_n6382 = n2716 & new_n6377;
  assign new_n6383 = n2715 & new_n6377;
  assign new_n6384 = n2714 & new_n6377;
  assign new_n6385 = n2713 & new_n6377;
  assign new_n6386 = new_n5500 & new_n6372;
  assign new_n6387 = ~new_n6386 & new_n6375;
  assign new_n6388 = n2712 & new_n6387;
  assign new_n6389 = n2711 & new_n6387;
  assign new_n6390 = n2710 & new_n6387;
  assign new_n6391 = n2709 & new_n6387;
  assign new_n6392 = n2708 & new_n6387;
  assign new_n6393 = n2707 & new_n6387;
  assign new_n6394 = n2706 & new_n6387;
  assign new_n6395 = n2705 & new_n6387;
  assign new_n6396 = new_n5433 & new_n6372;
  assign new_n6397 = ~new_n6374 & ~new_n6396;
  assign new_n6398 = new_n5513 & new_n6372;
  assign new_n6399 = ~new_n6398 & new_n6397;
  assign new_n6400 = n2704 & new_n6399;
  assign new_n6401 = n2703 & new_n6399;
  assign new_n6402 = n2702 & new_n6399;
  assign new_n6403 = n2701 & new_n6399;
  assign new_n6404 = n2700 & new_n6399;
  assign new_n6405 = n2699 & new_n6399;
  assign new_n6406 = n2698 & new_n6399;
  assign new_n6407 = n2697 & new_n6399;
  assign new_n6408 = new_n5524 & new_n6372;
  assign new_n6409 = ~new_n6408 & new_n6397;
  assign new_n6410 = n2696 & new_n6409;
  assign new_n6411 = n2695 & new_n6409;
  assign new_n6412 = n2694 & new_n6409;
  assign new_n6413 = n2693 & new_n6409;
  assign new_n6414 = n2692 & new_n6409;
  assign new_n6415 = n2691 & new_n6409;
  assign new_n6416 = n2690 & new_n6409;
  assign new_n6417 = n2689 & new_n6409;
  assign new_n6418 = new_n5484 & new_n6187;
  assign new_n6419 = new_n5434 & new_n6418;
  assign new_n6420 = new_n5430 & new_n6418;
  assign new_n6421 = ~new_n6419 & ~new_n6420;
  assign new_n6422 = new_n5438 & new_n6418;
  assign new_n6423 = ~new_n6422 & new_n6421;
  assign new_n6424 = n2752 & new_n6423;
  assign new_n6425 = n2751 & new_n6423;
  assign new_n6426 = n2750 & new_n6423;
  assign new_n6427 = n2749 & new_n6423;
  assign new_n6428 = n2748 & new_n6423;
  assign new_n6429 = n2747 & new_n6423;
  assign new_n6430 = n2746 & new_n6423;
  assign new_n6431 = n2745 & new_n6423;
  assign new_n6432 = new_n5500 & new_n6418;
  assign new_n6433 = ~new_n6432 & new_n6421;
  assign new_n6434 = n2744 & new_n6433;
  assign new_n6435 = n2743 & new_n6433;
  assign new_n6436 = n2742 & new_n6433;
  assign new_n6437 = n2741 & new_n6433;
  assign new_n6438 = n2740 & new_n6433;
  assign new_n6439 = n2739 & new_n6433;
  assign new_n6440 = n2738 & new_n6433;
  assign new_n6441 = n2737 & new_n6433;
  assign new_n6442 = new_n5433 & new_n6418;
  assign new_n6443 = ~new_n6420 & ~new_n6442;
  assign new_n6444 = new_n5513 & new_n6418;
  assign new_n6445 = ~new_n6444 & new_n6443;
  assign new_n6446 = n2736 & new_n6445;
  assign new_n6447 = n2735 & new_n6445;
  assign new_n6448 = n2734 & new_n6445;
  assign new_n6449 = n2733 & new_n6445;
  assign new_n6450 = n2732 & new_n6445;
  assign new_n6451 = n2731 & new_n6445;
  assign new_n6452 = n2730 & new_n6445;
  assign new_n6453 = n2729 & new_n6445;
  assign new_n6454 = new_n5524 & new_n6418;
  assign new_n6455 = ~new_n6454 & new_n6443;
  assign new_n6456 = n2728 & new_n6455;
  assign new_n6457 = n2727 & new_n6455;
  assign new_n6458 = n2726 & new_n6455;
  assign new_n6459 = n2725 & new_n6455;
  assign new_n6460 = n2724 & new_n6455;
  assign new_n6461 = n2723 & new_n6455;
  assign new_n6462 = n2722 & new_n6455;
  assign new_n6463 = n2721 & new_n6455;
  assign new_n6464 = new_n5536 & new_n6187;
  assign new_n6465 = new_n5434 & new_n6464;
  assign new_n6466 = new_n5430 & new_n6464;
  assign new_n6467 = ~new_n6465 & ~new_n6466;
  assign new_n6468 = new_n5438 & new_n6464;
  assign new_n6469 = ~new_n6468 & new_n6467;
  assign new_n6470 = n2784 & new_n6469;
  assign new_n6471 = n2783 & new_n6469;
  assign new_n6472 = n2782 & new_n6469;
  assign new_n6473 = n2781 & new_n6469;
  assign new_n6474 = n2780 & new_n6469;
  assign new_n6475 = n2779 & new_n6469;
  assign new_n6476 = n2778 & new_n6469;
  assign new_n6477 = n2777 & new_n6469;
  assign new_n6478 = new_n5500 & new_n6464;
  assign new_n6479 = ~new_n6478 & new_n6467;
  assign new_n6480 = n2776 & new_n6479;
  assign new_n6481 = n2775 & new_n6479;
  assign new_n6482 = n2774 & new_n6479;
  assign new_n6483 = n2773 & new_n6479;
  assign new_n6484 = n2772 & new_n6479;
  assign new_n6485 = n2771 & new_n6479;
  assign new_n6486 = n2770 & new_n6479;
  assign new_n6487 = n2769 & new_n6479;
  assign new_n6488 = new_n5433 & new_n6464;
  assign new_n6489 = ~new_n6466 & ~new_n6488;
  assign new_n6490 = new_n5513 & new_n6464;
  assign new_n6491 = ~new_n6490 & new_n6489;
  assign new_n6492 = n2768 & new_n6491;
  assign new_n6493 = n2767 & new_n6491;
  assign new_n6494 = n2766 & new_n6491;
  assign new_n6495 = n2765 & new_n6491;
  assign new_n6496 = n2764 & new_n6491;
  assign new_n6497 = n2763 & new_n6491;
  assign new_n6498 = n2762 & new_n6491;
  assign new_n6499 = n2761 & new_n6491;
  assign new_n6500 = new_n5524 & new_n6464;
  assign new_n6501 = ~new_n6500 & new_n6489;
  assign new_n6502 = n2760 & new_n6501;
  assign new_n6503 = n2759 & new_n6501;
  assign new_n6504 = n2758 & new_n6501;
  assign new_n6505 = n2757 & new_n6501;
  assign new_n6506 = n2756 & new_n6501;
  assign new_n6507 = n2755 & new_n6501;
  assign new_n6508 = n2754 & new_n6501;
  assign new_n6509 = n2753 & new_n6501;
  assign new_n6510 = new_n5246 & new_n6187;
  assign new_n6511 = new_n5434 & new_n6510;
  assign new_n6512 = new_n5430 & new_n6510;
  assign new_n6513 = ~new_n6511 & ~new_n6512;
  assign new_n6514 = new_n5438 & new_n6510;
  assign new_n6515 = ~new_n6514 & new_n6513;
  assign new_n6516 = n2816 & new_n6515;
  assign new_n6517 = n2815 & new_n6515;
  assign new_n6518 = n2814 & new_n6515;
  assign new_n6519 = n2813 & new_n6515;
  assign new_n6520 = n2812 & new_n6515;
  assign new_n6521 = n2811 & new_n6515;
  assign new_n6522 = n2810 & new_n6515;
  assign new_n6523 = n2809 & new_n6515;
  assign new_n6524 = new_n5500 & new_n6510;
  assign new_n6525 = ~new_n6524 & new_n6513;
  assign new_n6526 = n2808 & new_n6525;
  assign new_n6527 = n2807 & new_n6525;
  assign new_n6528 = n2806 & new_n6525;
  assign new_n6529 = n2805 & new_n6525;
  assign new_n6530 = n2804 & new_n6525;
  assign new_n6531 = n2803 & new_n6525;
  assign new_n6532 = n2802 & new_n6525;
  assign new_n6533 = n2801 & new_n6525;
  assign new_n6534 = new_n5433 & new_n6510;
  assign new_n6535 = ~new_n6512 & ~new_n6534;
  assign new_n6536 = new_n5513 & new_n6510;
  assign new_n6537 = ~new_n6536 & new_n6535;
  assign new_n6538 = n2800 & new_n6537;
  assign new_n6539 = n2799 & new_n6537;
  assign new_n6540 = n2798 & new_n6537;
  assign new_n6541 = n2797 & new_n6537;
  assign new_n6542 = n2796 & new_n6537;
  assign new_n6543 = n2795 & new_n6537;
  assign new_n6544 = n2794 & new_n6537;
  assign new_n6545 = n2793 & new_n6537;
  assign new_n6546 = new_n5524 & new_n6510;
  assign new_n6547 = ~new_n6546 & new_n6535;
  assign new_n6548 = n2792 & new_n6547;
  assign new_n6549 = n2791 & new_n6547;
  assign new_n6550 = n2790 & new_n6547;
  assign new_n6551 = n2789 & new_n6547;
  assign new_n6552 = n2788 & new_n6547;
  assign new_n6553 = n2787 & new_n6547;
  assign new_n6554 = n2786 & new_n6547;
  assign new_n6555 = n2785 & new_n6547;
  assign new_n6556 = new_n5011 & new_n5139;
  assign new_n6557 = new_n5031 & new_n6556;
  assign new_n6558 = new_n6557 ^ new_n6556;
  assign new_n6559 = new_n5424 & new_n6558;
  assign new_n6560 = new_n5434 & new_n6559;
  assign new_n6561 = new_n5430 & new_n6559;
  assign new_n6562 = ~new_n6560 & ~new_n6561;
  assign new_n6563 = new_n5438 & new_n6559;
  assign new_n6564 = ~new_n6563 & new_n6562;
  assign new_n6565 = n2848 & new_n6564;
  assign new_n6566 = n2847 & new_n6564;
  assign new_n6567 = n2846 & new_n6564;
  assign new_n6568 = n2845 & new_n6564;
  assign new_n6569 = n2844 & new_n6564;
  assign new_n6570 = n2843 & new_n6564;
  assign new_n6571 = n2842 & new_n6564;
  assign new_n6572 = n2841 & new_n6564;
  assign new_n6573 = new_n5500 & new_n6559;
  assign new_n6574 = ~new_n6573 & new_n6562;
  assign new_n6575 = n2840 & new_n6574;
  assign new_n6576 = n2839 & new_n6574;
  assign new_n6577 = n2838 & new_n6574;
  assign new_n6578 = n2837 & new_n6574;
  assign new_n6579 = n2836 & new_n6574;
  assign new_n6580 = n2835 & new_n6574;
  assign new_n6581 = n2834 & new_n6574;
  assign new_n6582 = n2833 & new_n6574;
  assign new_n6583 = new_n5433 & new_n6559;
  assign new_n6584 = ~new_n6561 & ~new_n6583;
  assign new_n6585 = new_n5513 & new_n6559;
  assign new_n6586 = ~new_n6585 & new_n6584;
  assign new_n6587 = n2832 & new_n6586;
  assign new_n6588 = n2831 & new_n6586;
  assign new_n6589 = n2830 & new_n6586;
  assign new_n6590 = n2829 & new_n6586;
  assign new_n6591 = n2828 & new_n6586;
  assign new_n6592 = n2827 & new_n6586;
  assign new_n6593 = n2826 & new_n6586;
  assign new_n6594 = n2825 & new_n6586;
  assign new_n6595 = new_n5524 & new_n6559;
  assign new_n6596 = ~new_n6595 & new_n6584;
  assign new_n6597 = n2824 & new_n6596;
  assign new_n6598 = n2823 & new_n6596;
  assign new_n6599 = n2822 & new_n6596;
  assign new_n6600 = n2821 & new_n6596;
  assign new_n6601 = n2820 & new_n6596;
  assign new_n6602 = n2819 & new_n6596;
  assign new_n6603 = n2818 & new_n6596;
  assign new_n6604 = n2817 & new_n6596;
  assign new_n6605 = new_n5485 & new_n6558;
  assign new_n6606 = new_n5434 & new_n6605;
  assign new_n6607 = new_n5430 & new_n6605;
  assign new_n6608 = ~new_n6606 & ~new_n6607;
  assign new_n6609 = new_n5438 & new_n6605;
  assign new_n6610 = ~new_n6609 & new_n6608;
  assign new_n6611 = n2880 & new_n6610;
  assign new_n6612 = n2879 & new_n6610;
  assign new_n6613 = n2878 & new_n6610;
  assign new_n6614 = n2877 & new_n6610;
  assign new_n6615 = n2876 & new_n6610;
  assign new_n6616 = n2875 & new_n6610;
  assign new_n6617 = n2874 & new_n6610;
  assign new_n6618 = n2873 & new_n6610;
  assign new_n6619 = new_n5500 & new_n6605;
  assign new_n6620 = ~new_n6619 & new_n6608;
  assign new_n6621 = n2872 & new_n6620;
  assign new_n6622 = n2871 & new_n6620;
  assign new_n6623 = n2870 & new_n6620;
  assign new_n6624 = n2869 & new_n6620;
  assign new_n6625 = n2868 & new_n6620;
  assign new_n6626 = n2867 & new_n6620;
  assign new_n6627 = n2866 & new_n6620;
  assign new_n6628 = n2865 & new_n6620;
  assign new_n6629 = new_n5433 & new_n6605;
  assign new_n6630 = ~new_n6607 & ~new_n6629;
  assign new_n6631 = new_n5513 & new_n6605;
  assign new_n6632 = ~new_n6631 & new_n6630;
  assign new_n6633 = n2864 & new_n6632;
  assign new_n6634 = n2863 & new_n6632;
  assign new_n6635 = n2862 & new_n6632;
  assign new_n6636 = n2861 & new_n6632;
  assign new_n6637 = n2860 & new_n6632;
  assign new_n6638 = n2859 & new_n6632;
  assign new_n6639 = n2858 & new_n6632;
  assign new_n6640 = n2857 & new_n6632;
  assign new_n6641 = new_n5524 & new_n6605;
  assign new_n6642 = ~new_n6641 & new_n6630;
  assign new_n6643 = n2856 & new_n6642;
  assign new_n6644 = n2855 & new_n6642;
  assign new_n6645 = n2854 & new_n6642;
  assign new_n6646 = n2853 & new_n6642;
  assign new_n6647 = n2852 & new_n6642;
  assign new_n6648 = n2851 & new_n6642;
  assign new_n6649 = n2850 & new_n6642;
  assign new_n6650 = n2849 & new_n6642;
  assign new_n6651 = new_n5537 & new_n6558;
  assign new_n6652 = new_n5434 & new_n6651;
  assign new_n6653 = new_n5430 & new_n6651;
  assign new_n6654 = ~new_n6652 & ~new_n6653;
  assign new_n6655 = new_n5438 & new_n6651;
  assign new_n6656 = ~new_n6655 & new_n6654;
  assign new_n6657 = n2912 & new_n6656;
  assign new_n6658 = n2911 & new_n6656;
  assign new_n6659 = n2910 & new_n6656;
  assign new_n6660 = n2909 & new_n6656;
  assign new_n6661 = n2908 & new_n6656;
  assign new_n6662 = n2907 & new_n6656;
  assign new_n6663 = n2906 & new_n6656;
  assign new_n6664 = n2905 & new_n6656;
  assign new_n6665 = new_n5500 & new_n6651;
  assign new_n6666 = ~new_n6665 & new_n6654;
  assign new_n6667 = n2904 & new_n6666;
  assign new_n6668 = n2903 & new_n6666;
  assign new_n6669 = n2902 & new_n6666;
  assign new_n6670 = n2901 & new_n6666;
  assign new_n6671 = n2900 & new_n6666;
  assign new_n6672 = n2899 & new_n6666;
  assign new_n6673 = n2898 & new_n6666;
  assign new_n6674 = n2897 & new_n6666;
  assign new_n6675 = new_n5433 & new_n6651;
  assign new_n6676 = ~new_n6653 & ~new_n6675;
  assign new_n6677 = new_n5513 & new_n6651;
  assign new_n6678 = ~new_n6677 & new_n6676;
  assign new_n6679 = n2896 & new_n6678;
  assign new_n6680 = n2895 & new_n6678;
  assign new_n6681 = n2894 & new_n6678;
  assign new_n6682 = n2893 & new_n6678;
  assign new_n6683 = n2892 & new_n6678;
  assign new_n6684 = n2891 & new_n6678;
  assign new_n6685 = n2890 & new_n6678;
  assign new_n6686 = n2889 & new_n6678;
  assign new_n6687 = new_n5524 & new_n6651;
  assign new_n6688 = ~new_n6687 & new_n6676;
  assign new_n6689 = n2888 & new_n6688;
  assign new_n6690 = n2887 & new_n6688;
  assign new_n6691 = n2886 & new_n6688;
  assign new_n6692 = n2885 & new_n6688;
  assign new_n6693 = n2884 & new_n6688;
  assign new_n6694 = n2883 & new_n6688;
  assign new_n6695 = n2882 & new_n6688;
  assign new_n6696 = n2881 & new_n6688;
  assign new_n6697 = new_n5245 & new_n6558;
  assign new_n6698 = new_n5434 & new_n6697;
  assign new_n6699 = new_n5430 & new_n6697;
  assign new_n6700 = ~new_n6698 & ~new_n6699;
  assign new_n6701 = new_n5438 & new_n6697;
  assign new_n6702 = ~new_n6701 & new_n6700;
  assign new_n6703 = n2944 & new_n6702;
  assign new_n6704 = n2943 & new_n6702;
  assign new_n6705 = n2942 & new_n6702;
  assign new_n6706 = n2941 & new_n6702;
  assign new_n6707 = n2940 & new_n6702;
  assign new_n6708 = n2939 & new_n6702;
  assign new_n6709 = n2938 & new_n6702;
  assign new_n6710 = n2937 & new_n6702;
  assign new_n6711 = new_n5500 & new_n6697;
  assign new_n6712 = ~new_n6711 & new_n6700;
  assign new_n6713 = n2936 & new_n6712;
  assign new_n6714 = n2935 & new_n6712;
  assign new_n6715 = n2934 & new_n6712;
  assign new_n6716 = n2933 & new_n6712;
  assign new_n6717 = n2932 & new_n6712;
  assign new_n6718 = n2931 & new_n6712;
  assign new_n6719 = n2930 & new_n6712;
  assign new_n6720 = n2929 & new_n6712;
  assign new_n6721 = new_n5433 & new_n6697;
  assign new_n6722 = ~new_n6699 & ~new_n6721;
  assign new_n6723 = new_n5513 & new_n6697;
  assign new_n6724 = ~new_n6723 & new_n6722;
  assign new_n6725 = n2928 & new_n6724;
  assign new_n6726 = n2927 & new_n6724;
  assign new_n6727 = n2926 & new_n6724;
  assign new_n6728 = n2925 & new_n6724;
  assign new_n6729 = n2924 & new_n6724;
  assign new_n6730 = n2923 & new_n6724;
  assign new_n6731 = n2922 & new_n6724;
  assign new_n6732 = n2921 & new_n6724;
  assign new_n6733 = new_n5524 & new_n6697;
  assign new_n6734 = ~new_n6733 & new_n6722;
  assign new_n6735 = n2920 & new_n6734;
  assign new_n6736 = n2919 & new_n6734;
  assign new_n6737 = n2918 & new_n6734;
  assign new_n6738 = n2917 & new_n6734;
  assign new_n6739 = n2916 & new_n6734;
  assign new_n6740 = n2915 & new_n6734;
  assign new_n6741 = n2914 & new_n6734;
  assign new_n6742 = n2913 & new_n6734;
  assign new_n6743 = new_n5423 & new_n6558;
  assign new_n6744 = new_n5434 & new_n6743;
  assign new_n6745 = new_n5430 & new_n6743;
  assign new_n6746 = ~new_n6744 & ~new_n6745;
  assign new_n6747 = new_n5438 & new_n6743;
  assign new_n6748 = ~new_n6747 & new_n6746;
  assign new_n6749 = n2976 & new_n6748;
  assign new_n6750 = n2975 & new_n6748;
  assign new_n6751 = n2974 & new_n6748;
  assign new_n6752 = n2973 & new_n6748;
  assign new_n6753 = n2972 & new_n6748;
  assign new_n6754 = n2971 & new_n6748;
  assign new_n6755 = n2970 & new_n6748;
  assign new_n6756 = n2969 & new_n6748;
  assign new_n6757 = new_n5500 & new_n6743;
  assign new_n6758 = ~new_n6757 & new_n6746;
  assign new_n6759 = n2968 & new_n6758;
  assign new_n6760 = n2967 & new_n6758;
  assign new_n6761 = n2966 & new_n6758;
  assign new_n6762 = n2965 & new_n6758;
  assign new_n6763 = n2964 & new_n6758;
  assign new_n6764 = n2963 & new_n6758;
  assign new_n6765 = n2962 & new_n6758;
  assign new_n6766 = n2961 & new_n6758;
  assign new_n6767 = new_n5433 & new_n6743;
  assign new_n6768 = ~new_n6745 & ~new_n6767;
  assign new_n6769 = new_n5513 & new_n6743;
  assign new_n6770 = ~new_n6769 & new_n6768;
  assign new_n6771 = n2960 & new_n6770;
  assign new_n6772 = n2959 & new_n6770;
  assign new_n6773 = n2958 & new_n6770;
  assign new_n6774 = n2957 & new_n6770;
  assign new_n6775 = n2956 & new_n6770;
  assign new_n6776 = n2955 & new_n6770;
  assign new_n6777 = n2954 & new_n6770;
  assign new_n6778 = n2953 & new_n6770;
  assign new_n6779 = new_n5524 & new_n6743;
  assign new_n6780 = ~new_n6779 & new_n6768;
  assign new_n6781 = n2952 & new_n6780;
  assign new_n6782 = n2951 & new_n6780;
  assign new_n6783 = n2950 & new_n6780;
  assign new_n6784 = n2949 & new_n6780;
  assign new_n6785 = n2948 & new_n6780;
  assign new_n6786 = n2947 & new_n6780;
  assign new_n6787 = n2946 & new_n6780;
  assign new_n6788 = n2945 & new_n6780;
  assign new_n6789 = new_n5484 & new_n6558;
  assign new_n6790 = new_n5434 & new_n6789;
  assign new_n6791 = new_n5430 & new_n6789;
  assign new_n6792 = ~new_n6790 & ~new_n6791;
  assign new_n6793 = new_n5438 & new_n6789;
  assign new_n6794 = ~new_n6793 & new_n6792;
  assign new_n6795 = n3008 & new_n6794;
  assign new_n6796 = n3007 & new_n6794;
  assign new_n6797 = n3006 & new_n6794;
  assign new_n6798 = n3005 & new_n6794;
  assign new_n6799 = n3004 & new_n6794;
  assign new_n6800 = n3003 & new_n6794;
  assign new_n6801 = n3002 & new_n6794;
  assign new_n6802 = n3001 & new_n6794;
  assign new_n6803 = new_n5500 & new_n6789;
  assign new_n6804 = ~new_n6803 & new_n6792;
  assign new_n6805 = n3000 & new_n6804;
  assign new_n6806 = n2999 & new_n6804;
  assign new_n6807 = n2998 & new_n6804;
  assign new_n6808 = n2997 & new_n6804;
  assign new_n6809 = n2996 & new_n6804;
  assign new_n6810 = n2995 & new_n6804;
  assign new_n6811 = n2994 & new_n6804;
  assign new_n6812 = n2993 & new_n6804;
  assign new_n6813 = new_n5433 & new_n6789;
  assign new_n6814 = ~new_n6791 & ~new_n6813;
  assign new_n6815 = new_n5513 & new_n6789;
  assign new_n6816 = ~new_n6815 & new_n6814;
  assign new_n6817 = n2992 & new_n6816;
  assign new_n6818 = n2991 & new_n6816;
  assign new_n6819 = n2990 & new_n6816;
  assign new_n6820 = n2989 & new_n6816;
  assign new_n6821 = n2988 & new_n6816;
  assign new_n6822 = n2987 & new_n6816;
  assign new_n6823 = n2986 & new_n6816;
  assign new_n6824 = n2985 & new_n6816;
  assign new_n6825 = new_n5524 & new_n6789;
  assign new_n6826 = ~new_n6825 & new_n6814;
  assign new_n6827 = n2984 & new_n6826;
  assign new_n6828 = n2983 & new_n6826;
  assign new_n6829 = n2982 & new_n6826;
  assign new_n6830 = n2981 & new_n6826;
  assign new_n6831 = n2980 & new_n6826;
  assign new_n6832 = n2979 & new_n6826;
  assign new_n6833 = n2978 & new_n6826;
  assign new_n6834 = n2977 & new_n6826;
  assign new_n6835 = new_n5536 & new_n6558;
  assign new_n6836 = new_n5434 & new_n6835;
  assign new_n6837 = new_n5430 & new_n6835;
  assign new_n6838 = ~new_n6836 & ~new_n6837;
  assign new_n6839 = new_n5438 & new_n6835;
  assign new_n6840 = ~new_n6839 & new_n6838;
  assign new_n6841 = n3040 & new_n6840;
  assign new_n6842 = n3039 & new_n6840;
  assign new_n6843 = n3038 & new_n6840;
  assign new_n6844 = n3037 & new_n6840;
  assign new_n6845 = n3036 & new_n6840;
  assign new_n6846 = n3035 & new_n6840;
  assign new_n6847 = n3034 & new_n6840;
  assign new_n6848 = n3033 & new_n6840;
  assign new_n6849 = new_n5500 & new_n6835;
  assign new_n6850 = ~new_n6849 & new_n6838;
  assign new_n6851 = n3032 & new_n6850;
  assign new_n6852 = n3031 & new_n6850;
  assign new_n6853 = n3030 & new_n6850;
  assign new_n6854 = n3029 & new_n6850;
  assign new_n6855 = n3028 & new_n6850;
  assign new_n6856 = n3027 & new_n6850;
  assign new_n6857 = n3026 & new_n6850;
  assign new_n6858 = n3025 & new_n6850;
  assign new_n6859 = new_n5433 & new_n6835;
  assign new_n6860 = ~new_n6837 & ~new_n6859;
  assign new_n6861 = new_n5513 & new_n6835;
  assign new_n6862 = ~new_n6861 & new_n6860;
  assign new_n6863 = n3024 & new_n6862;
  assign new_n6864 = n3023 & new_n6862;
  assign new_n6865 = n3022 & new_n6862;
  assign new_n6866 = n3021 & new_n6862;
  assign new_n6867 = n3020 & new_n6862;
  assign new_n6868 = n3019 & new_n6862;
  assign new_n6869 = n3018 & new_n6862;
  assign new_n6870 = n3017 & new_n6862;
  assign new_n6871 = new_n5524 & new_n6835;
  assign new_n6872 = ~new_n6871 & new_n6860;
  assign new_n6873 = n3016 & new_n6872;
  assign new_n6874 = n3015 & new_n6872;
  assign new_n6875 = n3014 & new_n6872;
  assign new_n6876 = n3013 & new_n6872;
  assign new_n6877 = n3012 & new_n6872;
  assign new_n6878 = n3011 & new_n6872;
  assign new_n6879 = n3010 & new_n6872;
  assign new_n6880 = n3009 & new_n6872;
  assign new_n6881 = new_n5246 & new_n6558;
  assign new_n6882 = new_n5434 & new_n6881;
  assign new_n6883 = new_n5430 & new_n6881;
  assign new_n6884 = ~new_n6882 & ~new_n6883;
  assign new_n6885 = new_n5438 & new_n6881;
  assign new_n6886 = ~new_n6885 & new_n6884;
  assign new_n6887 = n3072 & new_n6886;
  assign new_n6888 = n3071 & new_n6886;
  assign new_n6889 = n3070 & new_n6886;
  assign new_n6890 = n3069 & new_n6886;
  assign new_n6891 = n3068 & new_n6886;
  assign new_n6892 = n3067 & new_n6886;
  assign new_n6893 = n3066 & new_n6886;
  assign new_n6894 = n3065 & new_n6886;
  assign new_n6895 = new_n5500 & new_n6881;
  assign new_n6896 = ~new_n6895 & new_n6884;
  assign new_n6897 = n3064 & new_n6896;
  assign new_n6898 = n3063 & new_n6896;
  assign new_n6899 = n3062 & new_n6896;
  assign new_n6900 = n3061 & new_n6896;
  assign new_n6901 = n3060 & new_n6896;
  assign new_n6902 = n3059 & new_n6896;
  assign new_n6903 = n3058 & new_n6896;
  assign new_n6904 = n3057 & new_n6896;
  assign new_n6905 = new_n5433 & new_n6881;
  assign new_n6906 = ~new_n6883 & ~new_n6905;
  assign new_n6907 = new_n5513 & new_n6881;
  assign new_n6908 = ~new_n6907 & new_n6906;
  assign new_n6909 = n3056 & new_n6908;
  assign new_n6910 = n3055 & new_n6908;
  assign new_n6911 = n3054 & new_n6908;
  assign new_n6912 = n3053 & new_n6908;
  assign new_n6913 = n3052 & new_n6908;
  assign new_n6914 = n3051 & new_n6908;
  assign new_n6915 = n3050 & new_n6908;
  assign new_n6916 = n3049 & new_n6908;
  assign new_n6917 = new_n5524 & new_n6881;
  assign new_n6918 = ~new_n6917 & new_n6906;
  assign new_n6919 = n3048 & new_n6918;
  assign new_n6920 = n3047 & new_n6918;
  assign new_n6921 = n3046 & new_n6918;
  assign new_n6922 = n3045 & new_n6918;
  assign new_n6923 = n3044 & new_n6918;
  assign new_n6924 = n3043 & new_n6918;
  assign new_n6925 = n3042 & new_n6918;
  assign new_n6926 = n3041 & new_n6918;
  assign new_n6927 = new_n5424 & new_n5426;
  assign new_n6928 = new_n5434 & new_n6927;
  assign new_n6929 = new_n5430 & new_n6927;
  assign new_n6930 = ~new_n6928 & ~new_n6929;
  assign new_n6931 = new_n5438 & new_n6927;
  assign new_n6932 = ~new_n6931 & new_n6930;
  assign new_n6933 = n3104 & new_n6932;
  assign new_n6934 = n3103 & new_n6932;
  assign new_n6935 = n3102 & new_n6932;
  assign new_n6936 = n3101 & new_n6932;
  assign new_n6937 = n3100 & new_n6932;
  assign new_n6938 = n3099 & new_n6932;
  assign new_n6939 = n3098 & new_n6932;
  assign new_n6940 = n3097 & new_n6932;
  assign new_n6941 = new_n5500 & new_n6927;
  assign new_n6942 = ~new_n6941 & new_n6930;
  assign new_n6943 = n3096 & new_n6942;
  assign new_n6944 = n3095 & new_n6942;
  assign new_n6945 = n3094 & new_n6942;
  assign new_n6946 = n3093 & new_n6942;
  assign new_n6947 = n3092 & new_n6942;
  assign new_n6948 = n3091 & new_n6942;
  assign new_n6949 = n3090 & new_n6942;
  assign new_n6950 = n3089 & new_n6942;
  assign new_n6951 = new_n5433 & new_n6927;
  assign new_n6952 = ~new_n6929 & ~new_n6951;
  assign new_n6953 = new_n5513 & new_n6927;
  assign new_n6954 = ~new_n6953 & new_n6952;
  assign new_n6955 = n3088 & new_n6954;
  assign new_n6956 = n3087 & new_n6954;
  assign new_n6957 = n3086 & new_n6954;
  assign new_n6958 = n3085 & new_n6954;
  assign new_n6959 = n3084 & new_n6954;
  assign new_n6960 = n3083 & new_n6954;
  assign new_n6961 = n3082 & new_n6954;
  assign new_n6962 = n3081 & new_n6954;
  assign new_n6963 = new_n5524 & new_n6927;
  assign new_n6964 = ~new_n6963 & new_n6952;
  assign new_n6965 = n3080 & new_n6964;
  assign new_n6966 = n3079 & new_n6964;
  assign new_n6967 = n3078 & new_n6964;
  assign new_n6968 = n3077 & new_n6964;
  assign new_n6969 = n3076 & new_n6964;
  assign new_n6970 = n3075 & new_n6964;
  assign new_n6971 = n3074 & new_n6964;
  assign new_n6972 = n3073 & new_n6964;
  assign new_n6973 = new_n5426 & new_n5485;
  assign new_n6974 = new_n5434 & new_n6973;
  assign new_n6975 = new_n5430 & new_n6973;
  assign new_n6976 = ~new_n6974 & ~new_n6975;
  assign new_n6977 = new_n5438 & new_n6973;
  assign new_n6978 = ~new_n6977 & new_n6976;
  assign new_n6979 = n3136 & new_n6978;
  assign new_n6980 = n3135 & new_n6978;
  assign new_n6981 = n3134 & new_n6978;
  assign new_n6982 = n3133 & new_n6978;
  assign new_n6983 = n3132 & new_n6978;
  assign new_n6984 = n3131 & new_n6978;
  assign new_n6985 = n3130 & new_n6978;
  assign new_n6986 = n3129 & new_n6978;
  assign new_n6987 = new_n5500 & new_n6973;
  assign new_n6988 = ~new_n6987 & new_n6976;
  assign new_n6989 = n3128 & new_n6988;
  assign new_n6990 = n3127 & new_n6988;
  assign new_n6991 = n3126 & new_n6988;
  assign new_n6992 = n3125 & new_n6988;
  assign new_n6993 = n3124 & new_n6988;
  assign new_n6994 = n3123 & new_n6988;
  assign new_n6995 = n3122 & new_n6988;
  assign new_n6996 = n3121 & new_n6988;
  assign new_n6997 = new_n5433 & new_n6973;
  assign new_n6998 = ~new_n6975 & ~new_n6997;
  assign new_n6999 = new_n5513 & new_n6973;
  assign new_n7000 = ~new_n6999 & new_n6998;
  assign new_n7001 = n3120 & new_n7000;
  assign new_n7002 = n3119 & new_n7000;
  assign new_n7003 = n3118 & new_n7000;
  assign new_n7004 = n3117 & new_n7000;
  assign new_n7005 = n3116 & new_n7000;
  assign new_n7006 = n3115 & new_n7000;
  assign new_n7007 = n3114 & new_n7000;
  assign new_n7008 = n3113 & new_n7000;
  assign new_n7009 = new_n5524 & new_n6973;
  assign new_n7010 = ~new_n7009 & new_n6998;
  assign new_n7011 = n3112 & new_n7010;
  assign new_n7012 = n3111 & new_n7010;
  assign new_n7013 = n3110 & new_n7010;
  assign new_n7014 = n3109 & new_n7010;
  assign new_n7015 = n3108 & new_n7010;
  assign new_n7016 = n3107 & new_n7010;
  assign new_n7017 = n3106 & new_n7010;
  assign new_n7018 = n3105 & new_n7010;
  assign new_n7019 = new_n5426 & new_n5537;
  assign new_n7020 = new_n5434 & new_n7019;
  assign new_n7021 = new_n5430 & new_n7019;
  assign new_n7022 = ~new_n7020 & ~new_n7021;
  assign new_n7023 = new_n5438 & new_n7019;
  assign new_n7024 = ~new_n7023 & new_n7022;
  assign new_n7025 = n3168 & new_n7024;
  assign new_n7026 = n3167 & new_n7024;
  assign new_n7027 = n3166 & new_n7024;
  assign new_n7028 = n3165 & new_n7024;
  assign new_n7029 = n3164 & new_n7024;
  assign new_n7030 = n3163 & new_n7024;
  assign new_n7031 = n3162 & new_n7024;
  assign new_n7032 = n3161 & new_n7024;
  assign new_n7033 = new_n5500 & new_n7019;
  assign new_n7034 = ~new_n7033 & new_n7022;
  assign new_n7035 = n3160 & new_n7034;
  assign new_n7036 = n3159 & new_n7034;
  assign new_n7037 = n3158 & new_n7034;
  assign new_n7038 = n3157 & new_n7034;
  assign new_n7039 = n3156 & new_n7034;
  assign new_n7040 = n3155 & new_n7034;
  assign new_n7041 = n3154 & new_n7034;
  assign new_n7042 = n3153 & new_n7034;
  assign new_n7043 = new_n5433 & new_n7019;
  assign new_n7044 = ~new_n7021 & ~new_n7043;
  assign new_n7045 = new_n5513 & new_n7019;
  assign new_n7046 = ~new_n7045 & new_n7044;
  assign new_n7047 = n3152 & new_n7046;
  assign new_n7048 = n3151 & new_n7046;
  assign new_n7049 = n3150 & new_n7046;
  assign new_n7050 = n3149 & new_n7046;
  assign new_n7051 = n3148 & new_n7046;
  assign new_n7052 = n3147 & new_n7046;
  assign new_n7053 = n3146 & new_n7046;
  assign new_n7054 = n3145 & new_n7046;
  assign new_n7055 = new_n5524 & new_n7019;
  assign new_n7056 = ~new_n7055 & new_n7044;
  assign new_n7057 = n3144 & new_n7056;
  assign new_n7058 = n3143 & new_n7056;
  assign new_n7059 = n3142 & new_n7056;
  assign new_n7060 = n3141 & new_n7056;
  assign new_n7061 = n3140 & new_n7056;
  assign new_n7062 = n3139 & new_n7056;
  assign new_n7063 = n3138 & new_n7056;
  assign new_n7064 = n3137 & new_n7056;
  assign new_n7065 = new_n5245 & new_n5426;
  assign new_n7066 = new_n5434 & new_n7065;
  assign new_n7067 = new_n5430 & new_n7065;
  assign new_n7068 = ~new_n7066 & ~new_n7067;
  assign new_n7069 = new_n5438 & new_n7065;
  assign new_n7070 = ~new_n7069 & new_n7068;
  assign new_n7071 = n3200 & new_n7070;
  assign new_n7072 = n3199 & new_n7070;
  assign new_n7073 = n3198 & new_n7070;
  assign new_n7074 = n3197 & new_n7070;
  assign new_n7075 = n3196 & new_n7070;
  assign new_n7076 = n3195 & new_n7070;
  assign new_n7077 = n3194 & new_n7070;
  assign new_n7078 = n3193 & new_n7070;
  assign new_n7079 = new_n5500 & new_n7065;
  assign new_n7080 = ~new_n7079 & new_n7068;
  assign new_n7081 = n3192 & new_n7080;
  assign new_n7082 = n3191 & new_n7080;
  assign new_n7083 = n3190 & new_n7080;
  assign new_n7084 = n3189 & new_n7080;
  assign new_n7085 = n3188 & new_n7080;
  assign new_n7086 = n3187 & new_n7080;
  assign new_n7087 = n3186 & new_n7080;
  assign new_n7088 = n3185 & new_n7080;
  assign new_n7089 = new_n5433 & new_n7065;
  assign new_n7090 = ~new_n7067 & ~new_n7089;
  assign new_n7091 = new_n5513 & new_n7065;
  assign new_n7092 = ~new_n7091 & new_n7090;
  assign new_n7093 = n3184 & new_n7092;
  assign new_n7094 = n3183 & new_n7092;
  assign new_n7095 = n3182 & new_n7092;
  assign new_n7096 = n3181 & new_n7092;
  assign new_n7097 = n3180 & new_n7092;
  assign new_n7098 = n3179 & new_n7092;
  assign new_n7099 = n3178 & new_n7092;
  assign new_n7100 = n3177 & new_n7092;
  assign new_n7101 = new_n5524 & new_n7065;
  assign new_n7102 = ~new_n7101 & new_n7090;
  assign new_n7103 = n3176 & new_n7102;
  assign new_n7104 = n3175 & new_n7102;
  assign new_n7105 = n3174 & new_n7102;
  assign new_n7106 = n3173 & new_n7102;
  assign new_n7107 = n3172 & new_n7102;
  assign new_n7108 = n3171 & new_n7102;
  assign new_n7109 = n3170 & new_n7102;
  assign new_n7110 = n3169 & new_n7102;
  assign new_n7111 = new_n5423 & new_n5426;
  assign new_n7112 = new_n5434 & new_n7111;
  assign new_n7113 = new_n5430 & new_n7111;
  assign new_n7114 = ~new_n7112 & ~new_n7113;
  assign new_n7115 = new_n5438 & new_n7111;
  assign new_n7116 = ~new_n7115 & new_n7114;
  assign new_n7117 = n3232 & new_n7116;
  assign new_n7118 = n3231 & new_n7116;
  assign new_n7119 = n3230 & new_n7116;
  assign new_n7120 = n3229 & new_n7116;
  assign new_n7121 = n3228 & new_n7116;
  assign new_n7122 = n3227 & new_n7116;
  assign new_n7123 = n3226 & new_n7116;
  assign new_n7124 = n3225 & new_n7116;
  assign new_n7125 = new_n5500 & new_n7111;
  assign new_n7126 = ~new_n7125 & new_n7114;
  assign new_n7127 = n3224 & new_n7126;
  assign new_n7128 = n3223 & new_n7126;
  assign new_n7129 = n3222 & new_n7126;
  assign new_n7130 = n3221 & new_n7126;
  assign new_n7131 = n3220 & new_n7126;
  assign new_n7132 = n3219 & new_n7126;
  assign new_n7133 = n3218 & new_n7126;
  assign new_n7134 = n3217 & new_n7126;
  assign new_n7135 = new_n5433 & new_n7111;
  assign new_n7136 = ~new_n7113 & ~new_n7135;
  assign new_n7137 = new_n5513 & new_n7111;
  assign new_n7138 = ~new_n7137 & new_n7136;
  assign new_n7139 = n3216 & new_n7138;
  assign new_n7140 = n3215 & new_n7138;
  assign new_n7141 = n3214 & new_n7138;
  assign new_n7142 = n3213 & new_n7138;
  assign new_n7143 = n3212 & new_n7138;
  assign new_n7144 = n3211 & new_n7138;
  assign new_n7145 = n3210 & new_n7138;
  assign new_n7146 = n3209 & new_n7138;
  assign new_n7147 = new_n5524 & new_n7111;
  assign new_n7148 = ~new_n7147 & new_n7136;
  assign new_n7149 = n3208 & new_n7148;
  assign new_n7150 = n3207 & new_n7148;
  assign new_n7151 = n3206 & new_n7148;
  assign new_n7152 = n3205 & new_n7148;
  assign new_n7153 = n3204 & new_n7148;
  assign new_n7154 = n3203 & new_n7148;
  assign new_n7155 = n3202 & new_n7148;
  assign new_n7156 = n3201 & new_n7148;
  assign new_n7157 = new_n5426 & new_n5484;
  assign new_n7158 = new_n5434 & new_n7157;
  assign new_n7159 = new_n5430 & new_n7157;
  assign new_n7160 = ~new_n7158 & ~new_n7159;
  assign new_n7161 = new_n5438 & new_n7157;
  assign new_n7162 = ~new_n7161 & new_n7160;
  assign new_n7163 = n3264 & new_n7162;
  assign new_n7164 = n3263 & new_n7162;
  assign new_n7165 = n3262 & new_n7162;
  assign new_n7166 = n3261 & new_n7162;
  assign new_n7167 = n3260 & new_n7162;
  assign new_n7168 = n3259 & new_n7162;
  assign new_n7169 = n3258 & new_n7162;
  assign new_n7170 = n3257 & new_n7162;
  assign new_n7171 = new_n5500 & new_n7157;
  assign new_n7172 = ~new_n7171 & new_n7160;
  assign new_n7173 = n3256 & new_n7172;
  assign new_n7174 = n3255 & new_n7172;
  assign new_n7175 = n3254 & new_n7172;
  assign new_n7176 = n3253 & new_n7172;
  assign new_n7177 = n3252 & new_n7172;
  assign new_n7178 = n3251 & new_n7172;
  assign new_n7179 = n3250 & new_n7172;
  assign new_n7180 = n3249 & new_n7172;
  assign new_n7181 = new_n5433 & new_n7157;
  assign new_n7182 = ~new_n7159 & ~new_n7181;
  assign new_n7183 = new_n5513 & new_n7157;
  assign new_n7184 = ~new_n7183 & new_n7182;
  assign new_n7185 = n3248 & new_n7184;
  assign new_n7186 = n3247 & new_n7184;
  assign new_n7187 = n3246 & new_n7184;
  assign new_n7188 = n3245 & new_n7184;
  assign new_n7189 = n3244 & new_n7184;
  assign new_n7190 = n3243 & new_n7184;
  assign new_n7191 = n3242 & new_n7184;
  assign new_n7192 = n3241 & new_n7184;
  assign new_n7193 = new_n5524 & new_n7157;
  assign new_n7194 = ~new_n7193 & new_n7182;
  assign new_n7195 = n3240 & new_n7194;
  assign new_n7196 = n3239 & new_n7194;
  assign new_n7197 = n3238 & new_n7194;
  assign new_n7198 = n3237 & new_n7194;
  assign new_n7199 = n3236 & new_n7194;
  assign new_n7200 = n3235 & new_n7194;
  assign new_n7201 = n3234 & new_n7194;
  assign new_n7202 = n3233 & new_n7194;
  assign new_n7203 = new_n5426 & new_n5536;
  assign new_n7204 = new_n5434 & new_n7203;
  assign new_n7205 = new_n5430 & new_n7203;
  assign new_n7206 = ~new_n7204 & ~new_n7205;
  assign new_n7207 = new_n5438 & new_n7203;
  assign new_n7208 = ~new_n7207 & new_n7206;
  assign new_n7209 = n3296 & new_n7208;
  assign new_n7210 = n3295 & new_n7208;
  assign new_n7211 = n3294 & new_n7208;
  assign new_n7212 = n3293 & new_n7208;
  assign new_n7213 = n3292 & new_n7208;
  assign new_n7214 = n3291 & new_n7208;
  assign new_n7215 = n3290 & new_n7208;
  assign new_n7216 = n3289 & new_n7208;
  assign new_n7217 = new_n5500 & new_n7203;
  assign new_n7218 = ~new_n7217 & new_n7206;
  assign new_n7219 = n3288 & new_n7218;
  assign new_n7220 = n3287 & new_n7218;
  assign new_n7221 = n3286 & new_n7218;
  assign new_n7222 = n3285 & new_n7218;
  assign new_n7223 = n3284 & new_n7218;
  assign new_n7224 = n3283 & new_n7218;
  assign new_n7225 = n3282 & new_n7218;
  assign new_n7226 = n3281 & new_n7218;
  assign new_n7227 = new_n5433 & new_n7203;
  assign new_n7228 = ~new_n7205 & ~new_n7227;
  assign new_n7229 = new_n5513 & new_n7203;
  assign new_n7230 = ~new_n7229 & new_n7228;
  assign new_n7231 = n3280 & new_n7230;
  assign new_n7232 = n3279 & new_n7230;
  assign new_n7233 = n3278 & new_n7230;
  assign new_n7234 = n3277 & new_n7230;
  assign new_n7235 = n3276 & new_n7230;
  assign new_n7236 = n3275 & new_n7230;
  assign new_n7237 = n3274 & new_n7230;
  assign new_n7238 = n3273 & new_n7230;
  assign new_n7239 = new_n5524 & new_n7203;
  assign new_n7240 = ~new_n7239 & new_n7228;
  assign new_n7241 = n3272 & new_n7240;
  assign new_n7242 = n3271 & new_n7240;
  assign new_n7243 = n3270 & new_n7240;
  assign new_n7244 = n3269 & new_n7240;
  assign new_n7245 = n3268 & new_n7240;
  assign new_n7246 = n3267 & new_n7240;
  assign new_n7247 = n3266 & new_n7240;
  assign new_n7248 = n3265 & new_n7240;
  assign new_n7249 = new_n5246 & new_n5426;
  assign new_n7250 = new_n5434 & new_n7249;
  assign new_n7251 = new_n5430 & new_n7249;
  assign new_n7252 = ~new_n7250 & ~new_n7251;
  assign new_n7253 = new_n5438 & new_n7249;
  assign new_n7254 = ~new_n7253 & new_n7252;
  assign new_n7255 = n3328 & new_n7254;
  assign new_n7256 = n3327 & new_n7254;
  assign new_n7257 = n3326 & new_n7254;
  assign new_n7258 = n3325 & new_n7254;
  assign new_n7259 = n3324 & new_n7254;
  assign new_n7260 = n3323 & new_n7254;
  assign new_n7261 = n3322 & new_n7254;
  assign new_n7262 = n3321 & new_n7254;
  assign new_n7263 = new_n5500 & new_n7249;
  assign new_n7264 = ~new_n7263 & new_n7252;
  assign new_n7265 = n3320 & new_n7264;
  assign new_n7266 = n3319 & new_n7264;
  assign new_n7267 = n3318 & new_n7264;
  assign new_n7268 = n3317 & new_n7264;
  assign new_n7269 = n3316 & new_n7264;
  assign new_n7270 = n3315 & new_n7264;
  assign new_n7271 = n3314 & new_n7264;
  assign new_n7272 = n3313 & new_n7264;
  assign new_n7273 = new_n5433 & new_n7249;
  assign new_n7274 = ~new_n7251 & ~new_n7273;
  assign new_n7275 = new_n5513 & new_n7249;
  assign new_n7276 = ~new_n7275 & new_n7274;
  assign new_n7277 = n3312 & new_n7276;
  assign new_n7278 = n3311 & new_n7276;
  assign new_n7279 = n3310 & new_n7276;
  assign new_n7280 = n3309 & new_n7276;
  assign new_n7281 = n3308 & new_n7276;
  assign new_n7282 = n3307 & new_n7276;
  assign new_n7283 = n3306 & new_n7276;
  assign new_n7284 = n3305 & new_n7276;
  assign new_n7285 = new_n5524 & new_n7249;
  assign new_n7286 = ~new_n7285 & new_n7274;
  assign new_n7287 = n3304 & new_n7286;
  assign new_n7288 = n3303 & new_n7286;
  assign new_n7289 = n3302 & new_n7286;
  assign new_n7290 = n3301 & new_n7286;
  assign new_n7291 = n3300 & new_n7286;
  assign new_n7292 = n3299 & new_n7286;
  assign new_n7293 = n3298 & new_n7286;
  assign new_n7294 = n3297 & new_n7286;
  assign new_n7295 = new_n5424 & new_n5815;
  assign new_n7296 = new_n5434 & new_n7295;
  assign new_n7297 = new_n5430 & new_n7295;
  assign new_n7298 = ~new_n7296 & ~new_n7297;
  assign new_n7299 = new_n5438 & new_n7295;
  assign new_n7300 = ~new_n7299 & new_n7298;
  assign new_n7301 = n3360 & new_n7300;
  assign new_n7302 = n3359 & new_n7300;
  assign new_n7303 = n3358 & new_n7300;
  assign new_n7304 = n3357 & new_n7300;
  assign new_n7305 = n3356 & new_n7300;
  assign new_n7306 = n3355 & new_n7300;
  assign new_n7307 = n3354 & new_n7300;
  assign new_n7308 = n3353 & new_n7300;
  assign new_n7309 = new_n5500 & new_n7295;
  assign new_n7310 = ~new_n7309 & new_n7298;
  assign new_n7311 = n3352 & new_n7310;
  assign new_n7312 = n3351 & new_n7310;
  assign new_n7313 = n3350 & new_n7310;
  assign new_n7314 = n3349 & new_n7310;
  assign new_n7315 = n3348 & new_n7310;
  assign new_n7316 = n3347 & new_n7310;
  assign new_n7317 = n3346 & new_n7310;
  assign new_n7318 = n3345 & new_n7310;
  assign new_n7319 = new_n5433 & new_n7295;
  assign new_n7320 = ~new_n7297 & ~new_n7319;
  assign new_n7321 = new_n5513 & new_n7295;
  assign new_n7322 = ~new_n7321 & new_n7320;
  assign new_n7323 = n3344 & new_n7322;
  assign new_n7324 = n3343 & new_n7322;
  assign new_n7325 = n3342 & new_n7322;
  assign new_n7326 = n3341 & new_n7322;
  assign new_n7327 = n3340 & new_n7322;
  assign new_n7328 = n3339 & new_n7322;
  assign new_n7329 = n3338 & new_n7322;
  assign new_n7330 = n3337 & new_n7322;
  assign new_n7331 = new_n5524 & new_n7295;
  assign new_n7332 = ~new_n7331 & new_n7320;
  assign new_n7333 = n3336 & new_n7332;
  assign new_n7334 = n3335 & new_n7332;
  assign new_n7335 = n3334 & new_n7332;
  assign new_n7336 = n3333 & new_n7332;
  assign new_n7337 = n3332 & new_n7332;
  assign new_n7338 = n3331 & new_n7332;
  assign new_n7339 = n3330 & new_n7332;
  assign new_n7340 = n3329 & new_n7332;
  assign new_n7341 = new_n5485 & new_n5815;
  assign new_n7342 = new_n5434 & new_n7341;
  assign new_n7343 = new_n5430 & new_n7341;
  assign new_n7344 = ~new_n7342 & ~new_n7343;
  assign new_n7345 = new_n5438 & new_n7341;
  assign new_n7346 = ~new_n7345 & new_n7344;
  assign new_n7347 = n3392 & new_n7346;
  assign new_n7348 = n3391 & new_n7346;
  assign new_n7349 = n3390 & new_n7346;
  assign new_n7350 = n3389 & new_n7346;
  assign new_n7351 = n3388 & new_n7346;
  assign new_n7352 = n3387 & new_n7346;
  assign new_n7353 = n3386 & new_n7346;
  assign new_n7354 = n3385 & new_n7346;
  assign new_n7355 = new_n5500 & new_n7341;
  assign new_n7356 = ~new_n7355 & new_n7344;
  assign new_n7357 = n3384 & new_n7356;
  assign new_n7358 = n3383 & new_n7356;
  assign new_n7359 = n3382 & new_n7356;
  assign new_n7360 = n3381 & new_n7356;
  assign new_n7361 = n3380 & new_n7356;
  assign new_n7362 = n3379 & new_n7356;
  assign new_n7363 = n3378 & new_n7356;
  assign new_n7364 = n3377 & new_n7356;
  assign new_n7365 = new_n5433 & new_n7341;
  assign new_n7366 = ~new_n7343 & ~new_n7365;
  assign new_n7367 = new_n5513 & new_n7341;
  assign new_n7368 = ~new_n7367 & new_n7366;
  assign new_n7369 = n3376 & new_n7368;
  assign new_n7370 = n3375 & new_n7368;
  assign new_n7371 = n3374 & new_n7368;
  assign new_n7372 = n3373 & new_n7368;
  assign new_n7373 = n3372 & new_n7368;
  assign new_n7374 = n3371 & new_n7368;
  assign new_n7375 = n3370 & new_n7368;
  assign new_n7376 = n3369 & new_n7368;
  assign new_n7377 = new_n5524 & new_n7341;
  assign new_n7378 = ~new_n7377 & new_n7366;
  assign new_n7379 = n3368 & new_n7378;
  assign new_n7380 = n3367 & new_n7378;
  assign new_n7381 = n3366 & new_n7378;
  assign new_n7382 = n3365 & new_n7378;
  assign new_n7383 = n3364 & new_n7378;
  assign new_n7384 = n3363 & new_n7378;
  assign new_n7385 = n3362 & new_n7378;
  assign new_n7386 = n3361 & new_n7378;
  assign new_n7387 = new_n5537 & new_n5815;
  assign new_n7388 = new_n5434 & new_n7387;
  assign new_n7389 = new_n5430 & new_n7387;
  assign new_n7390 = ~new_n7388 & ~new_n7389;
  assign new_n7391 = new_n5438 & new_n7387;
  assign new_n7392 = ~new_n7391 & new_n7390;
  assign new_n7393 = n3424 & new_n7392;
  assign new_n7394 = n3423 & new_n7392;
  assign new_n7395 = n3422 & new_n7392;
  assign new_n7396 = n3421 & new_n7392;
  assign new_n7397 = n3420 & new_n7392;
  assign new_n7398 = n3419 & new_n7392;
  assign new_n7399 = n3418 & new_n7392;
  assign new_n7400 = n3417 & new_n7392;
  assign new_n7401 = new_n5500 & new_n7387;
  assign new_n7402 = ~new_n7401 & new_n7390;
  assign new_n7403 = n3416 & new_n7402;
  assign new_n7404 = n3415 & new_n7402;
  assign new_n7405 = n3414 & new_n7402;
  assign new_n7406 = n3413 & new_n7402;
  assign new_n7407 = n3412 & new_n7402;
  assign new_n7408 = n3411 & new_n7402;
  assign new_n7409 = n3410 & new_n7402;
  assign new_n7410 = n3409 & new_n7402;
  assign new_n7411 = new_n5433 & new_n7387;
  assign new_n7412 = ~new_n7389 & ~new_n7411;
  assign new_n7413 = new_n5513 & new_n7387;
  assign new_n7414 = ~new_n7413 & new_n7412;
  assign new_n7415 = n3408 & new_n7414;
  assign new_n7416 = n3407 & new_n7414;
  assign new_n7417 = n3406 & new_n7414;
  assign new_n7418 = n3405 & new_n7414;
  assign new_n7419 = n3404 & new_n7414;
  assign new_n7420 = n3403 & new_n7414;
  assign new_n7421 = n3402 & new_n7414;
  assign new_n7422 = n3401 & new_n7414;
  assign new_n7423 = new_n5524 & new_n7387;
  assign new_n7424 = ~new_n7423 & new_n7412;
  assign new_n7425 = n3400 & new_n7424;
  assign new_n7426 = n3399 & new_n7424;
  assign new_n7427 = n3398 & new_n7424;
  assign new_n7428 = n3397 & new_n7424;
  assign new_n7429 = n3396 & new_n7424;
  assign new_n7430 = n3395 & new_n7424;
  assign new_n7431 = n3394 & new_n7424;
  assign new_n7432 = n3393 & new_n7424;
  assign new_n7433 = new_n5245 & new_n5815;
  assign new_n7434 = new_n5434 & new_n7433;
  assign new_n7435 = new_n5430 & new_n7433;
  assign new_n7436 = ~new_n7434 & ~new_n7435;
  assign new_n7437 = new_n5438 & new_n7433;
  assign new_n7438 = ~new_n7437 & new_n7436;
  assign new_n7439 = n3456 & new_n7438;
  assign new_n7440 = n3455 & new_n7438;
  assign new_n7441 = n3454 & new_n7438;
  assign new_n7442 = n3453 & new_n7438;
  assign new_n7443 = n3452 & new_n7438;
  assign new_n7444 = n3451 & new_n7438;
  assign new_n7445 = n3450 & new_n7438;
  assign new_n7446 = n3449 & new_n7438;
  assign new_n7447 = new_n5500 & new_n7433;
  assign new_n7448 = ~new_n7447 & new_n7436;
  assign new_n7449 = n3448 & new_n7448;
  assign new_n7450 = n3447 & new_n7448;
  assign new_n7451 = n3446 & new_n7448;
  assign new_n7452 = n3445 & new_n7448;
  assign new_n7453 = n3444 & new_n7448;
  assign new_n7454 = n3443 & new_n7448;
  assign new_n7455 = n3442 & new_n7448;
  assign new_n7456 = n3441 & new_n7448;
  assign new_n7457 = new_n5433 & new_n7433;
  assign new_n7458 = ~new_n7435 & ~new_n7457;
  assign new_n7459 = new_n5513 & new_n7433;
  assign new_n7460 = ~new_n7459 & new_n7458;
  assign new_n7461 = n3440 & new_n7460;
  assign new_n7462 = n3439 & new_n7460;
  assign new_n7463 = n3438 & new_n7460;
  assign new_n7464 = n3437 & new_n7460;
  assign new_n7465 = n3436 & new_n7460;
  assign new_n7466 = n3435 & new_n7460;
  assign new_n7467 = n3434 & new_n7460;
  assign new_n7468 = n3433 & new_n7460;
  assign new_n7469 = new_n5524 & new_n7433;
  assign new_n7470 = ~new_n7469 & new_n7458;
  assign new_n7471 = n3432 & new_n7470;
  assign new_n7472 = n3431 & new_n7470;
  assign new_n7473 = n3430 & new_n7470;
  assign new_n7474 = n3429 & new_n7470;
  assign new_n7475 = n3428 & new_n7470;
  assign new_n7476 = n3427 & new_n7470;
  assign new_n7477 = n3426 & new_n7470;
  assign new_n7478 = n3425 & new_n7470;
  assign new_n7479 = new_n5423 & new_n5815;
  assign new_n7480 = new_n5434 & new_n7479;
  assign new_n7481 = new_n5430 & new_n7479;
  assign new_n7482 = ~new_n7480 & ~new_n7481;
  assign new_n7483 = new_n5438 & new_n7479;
  assign new_n7484 = ~new_n7483 & new_n7482;
  assign new_n7485 = n3488 & new_n7484;
  assign new_n7486 = n3487 & new_n7484;
  assign new_n7487 = n3486 & new_n7484;
  assign new_n7488 = n3485 & new_n7484;
  assign new_n7489 = n3484 & new_n7484;
  assign new_n7490 = n3483 & new_n7484;
  assign new_n7491 = n3482 & new_n7484;
  assign new_n7492 = n3481 & new_n7484;
  assign new_n7493 = new_n5500 & new_n7479;
  assign new_n7494 = ~new_n7493 & new_n7482;
  assign new_n7495 = n3480 & new_n7494;
  assign new_n7496 = n3479 & new_n7494;
  assign new_n7497 = n3478 & new_n7494;
  assign new_n7498 = n3477 & new_n7494;
  assign new_n7499 = n3476 & new_n7494;
  assign new_n7500 = n3475 & new_n7494;
  assign new_n7501 = n3474 & new_n7494;
  assign new_n7502 = n3473 & new_n7494;
  assign new_n7503 = new_n5433 & new_n7479;
  assign new_n7504 = ~new_n7481 & ~new_n7503;
  assign new_n7505 = new_n5513 & new_n7479;
  assign new_n7506 = ~new_n7505 & new_n7504;
  assign new_n7507 = n3472 & new_n7506;
  assign new_n7508 = n3471 & new_n7506;
  assign new_n7509 = n3470 & new_n7506;
  assign new_n7510 = n3469 & new_n7506;
  assign new_n7511 = n3468 & new_n7506;
  assign new_n7512 = n3467 & new_n7506;
  assign new_n7513 = n3466 & new_n7506;
  assign new_n7514 = n3465 & new_n7506;
  assign new_n7515 = new_n5524 & new_n7479;
  assign new_n7516 = ~new_n7515 & new_n7504;
  assign new_n7517 = n3464 & new_n7516;
  assign new_n7518 = n3463 & new_n7516;
  assign new_n7519 = n3462 & new_n7516;
  assign new_n7520 = n3461 & new_n7516;
  assign new_n7521 = n3460 & new_n7516;
  assign new_n7522 = n3459 & new_n7516;
  assign new_n7523 = n3458 & new_n7516;
  assign new_n7524 = n3457 & new_n7516;
  assign new_n7525 = new_n5484 & new_n5815;
  assign new_n7526 = new_n5434 & new_n7525;
  assign new_n7527 = new_n5430 & new_n7525;
  assign new_n7528 = ~new_n7526 & ~new_n7527;
  assign new_n7529 = new_n5438 & new_n7525;
  assign new_n7530 = ~new_n7529 & new_n7528;
  assign new_n7531 = n3520 & new_n7530;
  assign new_n7532 = n3519 & new_n7530;
  assign new_n7533 = n3518 & new_n7530;
  assign new_n7534 = n3517 & new_n7530;
  assign new_n7535 = n3516 & new_n7530;
  assign new_n7536 = n3515 & new_n7530;
  assign new_n7537 = n3514 & new_n7530;
  assign new_n7538 = n3513 & new_n7530;
  assign new_n7539 = new_n5500 & new_n7525;
  assign new_n7540 = ~new_n7539 & new_n7528;
  assign new_n7541 = n3512 & new_n7540;
  assign new_n7542 = n3511 & new_n7540;
  assign new_n7543 = n3510 & new_n7540;
  assign new_n7544 = n3509 & new_n7540;
  assign new_n7545 = n3508 & new_n7540;
  assign new_n7546 = n3507 & new_n7540;
  assign new_n7547 = n3506 & new_n7540;
  assign new_n7548 = n3505 & new_n7540;
  assign new_n7549 = new_n5433 & new_n7525;
  assign new_n7550 = ~new_n7527 & ~new_n7549;
  assign new_n7551 = new_n5513 & new_n7525;
  assign new_n7552 = ~new_n7551 & new_n7550;
  assign new_n7553 = n3504 & new_n7552;
  assign new_n7554 = n3503 & new_n7552;
  assign new_n7555 = n3502 & new_n7552;
  assign new_n7556 = n3501 & new_n7552;
  assign new_n7557 = n3500 & new_n7552;
  assign new_n7558 = n3499 & new_n7552;
  assign new_n7559 = n3498 & new_n7552;
  assign new_n7560 = n3497 & new_n7552;
  assign new_n7561 = new_n5524 & new_n7525;
  assign new_n7562 = ~new_n7561 & new_n7550;
  assign new_n7563 = n3496 & new_n7562;
  assign new_n7564 = n3495 & new_n7562;
  assign new_n7565 = n3494 & new_n7562;
  assign new_n7566 = n3493 & new_n7562;
  assign new_n7567 = n3492 & new_n7562;
  assign new_n7568 = n3491 & new_n7562;
  assign new_n7569 = n3490 & new_n7562;
  assign new_n7570 = n3489 & new_n7562;
  assign new_n7571 = new_n5536 & new_n5815;
  assign new_n7572 = new_n5434 & new_n7571;
  assign new_n7573 = new_n5430 & new_n7571;
  assign new_n7574 = ~new_n7572 & ~new_n7573;
  assign new_n7575 = new_n5438 & new_n7571;
  assign new_n7576 = ~new_n7575 & new_n7574;
  assign new_n7577 = n3552 & new_n7576;
  assign new_n7578 = n3551 & new_n7576;
  assign new_n7579 = n3550 & new_n7576;
  assign new_n7580 = n3549 & new_n7576;
  assign new_n7581 = n3548 & new_n7576;
  assign new_n7582 = n3547 & new_n7576;
  assign new_n7583 = n3546 & new_n7576;
  assign new_n7584 = n3545 & new_n7576;
  assign new_n7585 = new_n5500 & new_n7571;
  assign new_n7586 = ~new_n7585 & new_n7574;
  assign new_n7587 = n3544 & new_n7586;
  assign new_n7588 = n3543 & new_n7586;
  assign new_n7589 = n3542 & new_n7586;
  assign new_n7590 = n3541 & new_n7586;
  assign new_n7591 = n3540 & new_n7586;
  assign new_n7592 = n3539 & new_n7586;
  assign new_n7593 = n3538 & new_n7586;
  assign new_n7594 = n3537 & new_n7586;
  assign new_n7595 = new_n5433 & new_n7571;
  assign new_n7596 = ~new_n7573 & ~new_n7595;
  assign new_n7597 = new_n5513 & new_n7571;
  assign new_n7598 = ~new_n7597 & new_n7596;
  assign new_n7599 = n3536 & new_n7598;
  assign new_n7600 = n3535 & new_n7598;
  assign new_n7601 = n3534 & new_n7598;
  assign new_n7602 = n3533 & new_n7598;
  assign new_n7603 = n3532 & new_n7598;
  assign new_n7604 = n3531 & new_n7598;
  assign new_n7605 = n3530 & new_n7598;
  assign new_n7606 = n3529 & new_n7598;
  assign new_n7607 = new_n5524 & new_n7571;
  assign new_n7608 = ~new_n7607 & new_n7596;
  assign new_n7609 = n3528 & new_n7608;
  assign new_n7610 = n3527 & new_n7608;
  assign new_n7611 = n3526 & new_n7608;
  assign new_n7612 = n3525 & new_n7608;
  assign new_n7613 = n3524 & new_n7608;
  assign new_n7614 = n3523 & new_n7608;
  assign new_n7615 = n3522 & new_n7608;
  assign new_n7616 = n3521 & new_n7608;
  assign new_n7617 = new_n5246 & new_n5815;
  assign new_n7618 = new_n5434 & new_n7617;
  assign new_n7619 = new_n5430 & new_n7617;
  assign new_n7620 = ~new_n7618 & ~new_n7619;
  assign new_n7621 = new_n5438 & new_n7617;
  assign new_n7622 = ~new_n7621 & new_n7620;
  assign new_n7623 = n3584 & new_n7622;
  assign new_n7624 = n3583 & new_n7622;
  assign new_n7625 = n3582 & new_n7622;
  assign new_n7626 = n3581 & new_n7622;
  assign new_n7627 = n3580 & new_n7622;
  assign new_n7628 = n3579 & new_n7622;
  assign new_n7629 = n3578 & new_n7622;
  assign new_n7630 = n3577 & new_n7622;
  assign new_n7631 = new_n5500 & new_n7617;
  assign new_n7632 = ~new_n7631 & new_n7620;
  assign new_n7633 = n3576 & new_n7632;
  assign new_n7634 = n3575 & new_n7632;
  assign new_n7635 = n3574 & new_n7632;
  assign new_n7636 = n3573 & new_n7632;
  assign new_n7637 = n3572 & new_n7632;
  assign new_n7638 = n3571 & new_n7632;
  assign new_n7639 = n3570 & new_n7632;
  assign new_n7640 = n3569 & new_n7632;
  assign new_n7641 = new_n5433 & new_n7617;
  assign new_n7642 = ~new_n7619 & ~new_n7641;
  assign new_n7643 = new_n5513 & new_n7617;
  assign new_n7644 = ~new_n7643 & new_n7642;
  assign new_n7645 = n3568 & new_n7644;
  assign new_n7646 = n3567 & new_n7644;
  assign new_n7647 = n3566 & new_n7644;
  assign new_n7648 = n3565 & new_n7644;
  assign new_n7649 = n3564 & new_n7644;
  assign new_n7650 = n3563 & new_n7644;
  assign new_n7651 = n3562 & new_n7644;
  assign new_n7652 = n3561 & new_n7644;
  assign new_n7653 = new_n5524 & new_n7617;
  assign new_n7654 = ~new_n7653 & new_n7642;
  assign new_n7655 = n3560 & new_n7654;
  assign new_n7656 = n3559 & new_n7654;
  assign new_n7657 = n3558 & new_n7654;
  assign new_n7658 = n3557 & new_n7654;
  assign new_n7659 = n3556 & new_n7654;
  assign new_n7660 = n3555 & new_n7654;
  assign new_n7661 = n3554 & new_n7654;
  assign new_n7662 = n3553 & new_n7654;
  assign new_n7663 = new_n5424 & new_n6186;
  assign new_n7664 = new_n5434 & new_n7663;
  assign new_n7665 = new_n5430 & new_n7663;
  assign new_n7666 = ~new_n7664 & ~new_n7665;
  assign new_n7667 = new_n5438 & new_n7663;
  assign new_n7668 = ~new_n7667 & new_n7666;
  assign new_n7669 = n3616 & new_n7668;
  assign new_n7670 = n3615 & new_n7668;
  assign new_n7671 = n3614 & new_n7668;
  assign new_n7672 = n3613 & new_n7668;
  assign new_n7673 = n3612 & new_n7668;
  assign new_n7674 = n3611 & new_n7668;
  assign new_n7675 = n3610 & new_n7668;
  assign new_n7676 = n3609 & new_n7668;
  assign new_n7677 = new_n5500 & new_n7663;
  assign new_n7678 = ~new_n7677 & new_n7666;
  assign new_n7679 = n3608 & new_n7678;
  assign new_n7680 = n3607 & new_n7678;
  assign new_n7681 = n3606 & new_n7678;
  assign new_n7682 = n3605 & new_n7678;
  assign new_n7683 = n3604 & new_n7678;
  assign new_n7684 = n3603 & new_n7678;
  assign new_n7685 = n3602 & new_n7678;
  assign new_n7686 = n3601 & new_n7678;
  assign new_n7687 = new_n5433 & new_n7663;
  assign new_n7688 = ~new_n7665 & ~new_n7687;
  assign new_n7689 = new_n5513 & new_n7663;
  assign new_n7690 = ~new_n7689 & new_n7688;
  assign new_n7691 = n3600 & new_n7690;
  assign new_n7692 = n3599 & new_n7690;
  assign new_n7693 = n3598 & new_n7690;
  assign new_n7694 = n3597 & new_n7690;
  assign new_n7695 = n3596 & new_n7690;
  assign new_n7696 = n3595 & new_n7690;
  assign new_n7697 = n3594 & new_n7690;
  assign new_n7698 = n3593 & new_n7690;
  assign new_n7699 = new_n5524 & new_n7663;
  assign new_n7700 = ~new_n7699 & new_n7688;
  assign new_n7701 = n3592 & new_n7700;
  assign new_n7702 = n3591 & new_n7700;
  assign new_n7703 = n3590 & new_n7700;
  assign new_n7704 = n3589 & new_n7700;
  assign new_n7705 = n3588 & new_n7700;
  assign new_n7706 = n3587 & new_n7700;
  assign new_n7707 = n3586 & new_n7700;
  assign new_n7708 = n3585 & new_n7700;
  assign new_n7709 = new_n5485 & new_n6186;
  assign new_n7710 = new_n5434 & new_n7709;
  assign new_n7711 = new_n5430 & new_n7709;
  assign new_n7712 = ~new_n7710 & ~new_n7711;
  assign new_n7713 = new_n5438 & new_n7709;
  assign new_n7714 = ~new_n7713 & new_n7712;
  assign new_n7715 = n3648 & new_n7714;
  assign new_n7716 = n3647 & new_n7714;
  assign new_n7717 = n3646 & new_n7714;
  assign new_n7718 = n3645 & new_n7714;
  assign new_n7719 = n3644 & new_n7714;
  assign new_n7720 = n3643 & new_n7714;
  assign new_n7721 = n3642 & new_n7714;
  assign new_n7722 = n3641 & new_n7714;
  assign new_n7723 = new_n5500 & new_n7709;
  assign new_n7724 = ~new_n7723 & new_n7712;
  assign new_n7725 = n3640 & new_n7724;
  assign new_n7726 = n3639 & new_n7724;
  assign new_n7727 = n3638 & new_n7724;
  assign new_n7728 = n3637 & new_n7724;
  assign new_n7729 = n3636 & new_n7724;
  assign new_n7730 = n3635 & new_n7724;
  assign new_n7731 = n3634 & new_n7724;
  assign new_n7732 = n3633 & new_n7724;
  assign new_n7733 = new_n5433 & new_n7709;
  assign new_n7734 = ~new_n7711 & ~new_n7733;
  assign new_n7735 = new_n5513 & new_n7709;
  assign new_n7736 = ~new_n7735 & new_n7734;
  assign new_n7737 = n3632 & new_n7736;
  assign new_n7738 = n3631 & new_n7736;
  assign new_n7739 = n3630 & new_n7736;
  assign new_n7740 = n3629 & new_n7736;
  assign new_n7741 = n3628 & new_n7736;
  assign new_n7742 = n3627 & new_n7736;
  assign new_n7743 = n3626 & new_n7736;
  assign new_n7744 = n3625 & new_n7736;
  assign new_n7745 = new_n5524 & new_n7709;
  assign new_n7746 = ~new_n7745 & new_n7734;
  assign new_n7747 = n3624 & new_n7746;
  assign new_n7748 = n3623 & new_n7746;
  assign new_n7749 = n3622 & new_n7746;
  assign new_n7750 = n3621 & new_n7746;
  assign new_n7751 = n3620 & new_n7746;
  assign new_n7752 = n3619 & new_n7746;
  assign new_n7753 = n3618 & new_n7746;
  assign new_n7754 = n3617 & new_n7746;
  assign new_n7755 = new_n5537 & new_n6186;
  assign new_n7756 = new_n5434 & new_n7755;
  assign new_n7757 = new_n5430 & new_n7755;
  assign new_n7758 = ~new_n7756 & ~new_n7757;
  assign new_n7759 = new_n5438 & new_n7755;
  assign new_n7760 = ~new_n7759 & new_n7758;
  assign new_n7761 = n3680 & new_n7760;
  assign new_n7762 = n3679 & new_n7760;
  assign new_n7763 = n3678 & new_n7760;
  assign new_n7764 = n3677 & new_n7760;
  assign new_n7765 = n3676 & new_n7760;
  assign new_n7766 = n3675 & new_n7760;
  assign new_n7767 = n3674 & new_n7760;
  assign new_n7768 = n3673 & new_n7760;
  assign new_n7769 = new_n5500 & new_n7755;
  assign new_n7770 = ~new_n7769 & new_n7758;
  assign new_n7771 = n3672 & new_n7770;
  assign new_n7772 = n3671 & new_n7770;
  assign new_n7773 = n3670 & new_n7770;
  assign new_n7774 = n3669 & new_n7770;
  assign new_n7775 = n3668 & new_n7770;
  assign new_n7776 = n3667 & new_n7770;
  assign new_n7777 = n3666 & new_n7770;
  assign new_n7778 = n3665 & new_n7770;
  assign new_n7779 = new_n5433 & new_n7755;
  assign new_n7780 = ~new_n7757 & ~new_n7779;
  assign new_n7781 = new_n5513 & new_n7755;
  assign new_n7782 = ~new_n7781 & new_n7780;
  assign new_n7783 = n3664 & new_n7782;
  assign new_n7784 = n3663 & new_n7782;
  assign new_n7785 = n3662 & new_n7782;
  assign new_n7786 = n3661 & new_n7782;
  assign new_n7787 = n3660 & new_n7782;
  assign new_n7788 = n3659 & new_n7782;
  assign new_n7789 = n3658 & new_n7782;
  assign new_n7790 = n3657 & new_n7782;
  assign new_n7791 = new_n5524 & new_n7755;
  assign new_n7792 = ~new_n7791 & new_n7780;
  assign new_n7793 = n3656 & new_n7792;
  assign new_n7794 = n3655 & new_n7792;
  assign new_n7795 = n3654 & new_n7792;
  assign new_n7796 = n3653 & new_n7792;
  assign new_n7797 = n3652 & new_n7792;
  assign new_n7798 = n3651 & new_n7792;
  assign new_n7799 = n3650 & new_n7792;
  assign new_n7800 = n3649 & new_n7792;
  assign new_n7801 = new_n5245 & new_n6186;
  assign new_n7802 = new_n5434 & new_n7801;
  assign new_n7803 = new_n5430 & new_n7801;
  assign new_n7804 = ~new_n7802 & ~new_n7803;
  assign new_n7805 = new_n5438 & new_n7801;
  assign new_n7806 = ~new_n7805 & new_n7804;
  assign new_n7807 = n3712 & new_n7806;
  assign new_n7808 = n3711 & new_n7806;
  assign new_n7809 = n3710 & new_n7806;
  assign new_n7810 = n3709 & new_n7806;
  assign new_n7811 = n3708 & new_n7806;
  assign new_n7812 = n3707 & new_n7806;
  assign new_n7813 = n3706 & new_n7806;
  assign new_n7814 = n3705 & new_n7806;
  assign new_n7815 = new_n5500 & new_n7801;
  assign new_n7816 = ~new_n7815 & new_n7804;
  assign new_n7817 = n3704 & new_n7816;
  assign new_n7818 = n3703 & new_n7816;
  assign new_n7819 = n3702 & new_n7816;
  assign new_n7820 = n3701 & new_n7816;
  assign new_n7821 = n3700 & new_n7816;
  assign new_n7822 = n3699 & new_n7816;
  assign new_n7823 = n3698 & new_n7816;
  assign new_n7824 = n3697 & new_n7816;
  assign new_n7825 = new_n5433 & new_n7801;
  assign new_n7826 = ~new_n7803 & ~new_n7825;
  assign new_n7827 = new_n5513 & new_n7801;
  assign new_n7828 = ~new_n7827 & new_n7826;
  assign new_n7829 = n3696 & new_n7828;
  assign new_n7830 = n3695 & new_n7828;
  assign new_n7831 = n3694 & new_n7828;
  assign new_n7832 = n3693 & new_n7828;
  assign new_n7833 = n3692 & new_n7828;
  assign new_n7834 = n3691 & new_n7828;
  assign new_n7835 = n3690 & new_n7828;
  assign new_n7836 = n3689 & new_n7828;
  assign new_n7837 = new_n5524 & new_n7801;
  assign new_n7838 = ~new_n7837 & new_n7826;
  assign new_n7839 = n3688 & new_n7838;
  assign new_n7840 = n3687 & new_n7838;
  assign new_n7841 = n3686 & new_n7838;
  assign new_n7842 = n3685 & new_n7838;
  assign new_n7843 = n3684 & new_n7838;
  assign new_n7844 = n3683 & new_n7838;
  assign new_n7845 = n3682 & new_n7838;
  assign new_n7846 = n3681 & new_n7838;
  assign new_n7847 = new_n5423 & new_n6186;
  assign new_n7848 = new_n5434 & new_n7847;
  assign new_n7849 = new_n5430 & new_n7847;
  assign new_n7850 = ~new_n7848 & ~new_n7849;
  assign new_n7851 = new_n5438 & new_n7847;
  assign new_n7852 = ~new_n7851 & new_n7850;
  assign new_n7853 = n3744 & new_n7852;
  assign new_n7854 = n3743 & new_n7852;
  assign new_n7855 = n3742 & new_n7852;
  assign new_n7856 = n3741 & new_n7852;
  assign new_n7857 = n3740 & new_n7852;
  assign new_n7858 = n3739 & new_n7852;
  assign new_n7859 = n3738 & new_n7852;
  assign new_n7860 = n3737 & new_n7852;
  assign new_n7861 = new_n5500 & new_n7847;
  assign new_n7862 = ~new_n7861 & new_n7850;
  assign new_n7863 = n3736 & new_n7862;
  assign new_n7864 = n3735 & new_n7862;
  assign new_n7865 = n3734 & new_n7862;
  assign new_n7866 = n3733 & new_n7862;
  assign new_n7867 = n3732 & new_n7862;
  assign new_n7868 = n3731 & new_n7862;
  assign new_n7869 = n3730 & new_n7862;
  assign new_n7870 = n3729 & new_n7862;
  assign new_n7871 = new_n5433 & new_n7847;
  assign new_n7872 = ~new_n7849 & ~new_n7871;
  assign new_n7873 = new_n5513 & new_n7847;
  assign new_n7874 = ~new_n7873 & new_n7872;
  assign new_n7875 = n3728 & new_n7874;
  assign new_n7876 = n3727 & new_n7874;
  assign new_n7877 = n3726 & new_n7874;
  assign new_n7878 = n3725 & new_n7874;
  assign new_n7879 = n3724 & new_n7874;
  assign new_n7880 = n3723 & new_n7874;
  assign new_n7881 = n3722 & new_n7874;
  assign new_n7882 = n3721 & new_n7874;
  assign new_n7883 = new_n5524 & new_n7847;
  assign new_n7884 = ~new_n7883 & new_n7872;
  assign new_n7885 = n3720 & new_n7884;
  assign new_n7886 = n3719 & new_n7884;
  assign new_n7887 = n3718 & new_n7884;
  assign new_n7888 = n3717 & new_n7884;
  assign new_n7889 = n3716 & new_n7884;
  assign new_n7890 = n3715 & new_n7884;
  assign new_n7891 = n3714 & new_n7884;
  assign new_n7892 = n3713 & new_n7884;
  assign new_n7893 = new_n5484 & new_n6186;
  assign new_n7894 = new_n5434 & new_n7893;
  assign new_n7895 = new_n5430 & new_n7893;
  assign new_n7896 = ~new_n7894 & ~new_n7895;
  assign new_n7897 = new_n5438 & new_n7893;
  assign new_n7898 = ~new_n7897 & new_n7896;
  assign new_n7899 = n3776 & new_n7898;
  assign new_n7900 = n3775 & new_n7898;
  assign new_n7901 = n3774 & new_n7898;
  assign new_n7902 = n3773 & new_n7898;
  assign new_n7903 = n3772 & new_n7898;
  assign new_n7904 = n3771 & new_n7898;
  assign new_n7905 = n3770 & new_n7898;
  assign new_n7906 = n3769 & new_n7898;
  assign new_n7907 = new_n5500 & new_n7893;
  assign new_n7908 = ~new_n7907 & new_n7896;
  assign new_n7909 = n3768 & new_n7908;
  assign new_n7910 = n3767 & new_n7908;
  assign new_n7911 = n3766 & new_n7908;
  assign new_n7912 = n3765 & new_n7908;
  assign new_n7913 = n3764 & new_n7908;
  assign new_n7914 = n3763 & new_n7908;
  assign new_n7915 = n3762 & new_n7908;
  assign new_n7916 = n3761 & new_n7908;
  assign new_n7917 = new_n5433 & new_n7893;
  assign new_n7918 = ~new_n7895 & ~new_n7917;
  assign new_n7919 = new_n5513 & new_n7893;
  assign new_n7920 = ~new_n7919 & new_n7918;
  assign new_n7921 = n3760 & new_n7920;
  assign new_n7922 = n3759 & new_n7920;
  assign new_n7923 = n3758 & new_n7920;
  assign new_n7924 = n3757 & new_n7920;
  assign new_n7925 = n3756 & new_n7920;
  assign new_n7926 = n3755 & new_n7920;
  assign new_n7927 = n3754 & new_n7920;
  assign new_n7928 = n3753 & new_n7920;
  assign new_n7929 = new_n5524 & new_n7893;
  assign new_n7930 = ~new_n7929 & new_n7918;
  assign new_n7931 = n3752 & new_n7930;
  assign new_n7932 = n3751 & new_n7930;
  assign new_n7933 = n3750 & new_n7930;
  assign new_n7934 = n3749 & new_n7930;
  assign new_n7935 = n3748 & new_n7930;
  assign new_n7936 = n3747 & new_n7930;
  assign new_n7937 = n3746 & new_n7930;
  assign new_n7938 = n3745 & new_n7930;
  assign new_n7939 = new_n5536 & new_n6186;
  assign new_n7940 = new_n5434 & new_n7939;
  assign new_n7941 = new_n5430 & new_n7939;
  assign new_n7942 = ~new_n7940 & ~new_n7941;
  assign new_n7943 = new_n5438 & new_n7939;
  assign new_n7944 = ~new_n7943 & new_n7942;
  assign new_n7945 = n3808 & new_n7944;
  assign new_n7946 = n3807 & new_n7944;
  assign new_n7947 = n3806 & new_n7944;
  assign new_n7948 = n3805 & new_n7944;
  assign new_n7949 = n3804 & new_n7944;
  assign new_n7950 = n3803 & new_n7944;
  assign new_n7951 = n3802 & new_n7944;
  assign new_n7952 = n3801 & new_n7944;
  assign new_n7953 = new_n5500 & new_n7939;
  assign new_n7954 = ~new_n7953 & new_n7942;
  assign new_n7955 = n3800 & new_n7954;
  assign new_n7956 = n3799 & new_n7954;
  assign new_n7957 = n3798 & new_n7954;
  assign new_n7958 = n3797 & new_n7954;
  assign new_n7959 = n3796 & new_n7954;
  assign new_n7960 = n3795 & new_n7954;
  assign new_n7961 = n3794 & new_n7954;
  assign new_n7962 = n3793 & new_n7954;
  assign new_n7963 = new_n5433 & new_n7939;
  assign new_n7964 = ~new_n7941 & ~new_n7963;
  assign new_n7965 = new_n5513 & new_n7939;
  assign new_n7966 = ~new_n7965 & new_n7964;
  assign new_n7967 = n3792 & new_n7966;
  assign new_n7968 = n3791 & new_n7966;
  assign new_n7969 = n3790 & new_n7966;
  assign new_n7970 = n3789 & new_n7966;
  assign new_n7971 = n3788 & new_n7966;
  assign new_n7972 = n3787 & new_n7966;
  assign new_n7973 = n3786 & new_n7966;
  assign new_n7974 = n3785 & new_n7966;
  assign new_n7975 = new_n5524 & new_n7939;
  assign new_n7976 = ~new_n7975 & new_n7964;
  assign new_n7977 = n3784 & new_n7976;
  assign new_n7978 = n3783 & new_n7976;
  assign new_n7979 = n3782 & new_n7976;
  assign new_n7980 = n3781 & new_n7976;
  assign new_n7981 = n3780 & new_n7976;
  assign new_n7982 = n3779 & new_n7976;
  assign new_n7983 = n3778 & new_n7976;
  assign new_n7984 = n3777 & new_n7976;
  assign new_n7985 = new_n5246 & new_n6186;
  assign new_n7986 = new_n5434 & new_n7985;
  assign new_n7987 = new_n5430 & new_n7985;
  assign new_n7988 = ~new_n7986 & ~new_n7987;
  assign new_n7989 = new_n5438 & new_n7985;
  assign new_n7990 = ~new_n7989 & new_n7988;
  assign new_n7991 = n3840 & new_n7990;
  assign new_n7992 = n3839 & new_n7990;
  assign new_n7993 = n3838 & new_n7990;
  assign new_n7994 = n3837 & new_n7990;
  assign new_n7995 = n3836 & new_n7990;
  assign new_n7996 = n3835 & new_n7990;
  assign new_n7997 = n3834 & new_n7990;
  assign new_n7998 = n3833 & new_n7990;
  assign new_n7999 = new_n5500 & new_n7985;
  assign new_n8000 = ~new_n7999 & new_n7988;
  assign new_n8001 = n3832 & new_n8000;
  assign new_n8002 = n3831 & new_n8000;
  assign new_n8003 = n3830 & new_n8000;
  assign new_n8004 = n3829 & new_n8000;
  assign new_n8005 = n3828 & new_n8000;
  assign new_n8006 = n3827 & new_n8000;
  assign new_n8007 = n3826 & new_n8000;
  assign new_n8008 = n3825 & new_n8000;
  assign new_n8009 = new_n5433 & new_n7985;
  assign new_n8010 = ~new_n7987 & ~new_n8009;
  assign new_n8011 = new_n5513 & new_n7985;
  assign new_n8012 = ~new_n8011 & new_n8010;
  assign new_n8013 = n3824 & new_n8012;
  assign new_n8014 = n3823 & new_n8012;
  assign new_n8015 = n3822 & new_n8012;
  assign new_n8016 = n3821 & new_n8012;
  assign new_n8017 = n3820 & new_n8012;
  assign new_n8018 = n3819 & new_n8012;
  assign new_n8019 = n3818 & new_n8012;
  assign new_n8020 = n3817 & new_n8012;
  assign new_n8021 = new_n5524 & new_n7985;
  assign new_n8022 = ~new_n8021 & new_n8010;
  assign new_n8023 = n3816 & new_n8022;
  assign new_n8024 = n3815 & new_n8022;
  assign new_n8025 = n3814 & new_n8022;
  assign new_n8026 = n3813 & new_n8022;
  assign new_n8027 = n3812 & new_n8022;
  assign new_n8028 = n3811 & new_n8022;
  assign new_n8029 = n3810 & new_n8022;
  assign new_n8030 = n3809 & new_n8022;
  assign new_n8031 = new_n5424 & new_n6557;
  assign new_n8032 = new_n5434 & new_n8031;
  assign new_n8033 = new_n5430 & new_n8031;
  assign new_n8034 = ~new_n8032 & ~new_n8033;
  assign new_n8035 = new_n5438 & new_n8031;
  assign new_n8036 = ~new_n8035 & new_n8034;
  assign new_n8037 = n3872 & new_n8036;
  assign new_n8038 = n3871 & new_n8036;
  assign new_n8039 = n3870 & new_n8036;
  assign new_n8040 = n3869 & new_n8036;
  assign new_n8041 = n3868 & new_n8036;
  assign new_n8042 = n3867 & new_n8036;
  assign new_n8043 = n3866 & new_n8036;
  assign new_n8044 = n3865 & new_n8036;
  assign new_n8045 = new_n5500 & new_n8031;
  assign new_n8046 = ~new_n8045 & new_n8034;
  assign new_n8047 = n3864 & new_n8046;
  assign new_n8048 = n3863 & new_n8046;
  assign new_n8049 = n3862 & new_n8046;
  assign new_n8050 = n3861 & new_n8046;
  assign new_n8051 = n3860 & new_n8046;
  assign new_n8052 = n3859 & new_n8046;
  assign new_n8053 = n3858 & new_n8046;
  assign new_n8054 = n3857 & new_n8046;
  assign new_n8055 = new_n5433 & new_n8031;
  assign new_n8056 = ~new_n8033 & ~new_n8055;
  assign new_n8057 = new_n5513 & new_n8031;
  assign new_n8058 = ~new_n8057 & new_n8056;
  assign new_n8059 = n3856 & new_n8058;
  assign new_n8060 = n3855 & new_n8058;
  assign new_n8061 = n3854 & new_n8058;
  assign new_n8062 = n3853 & new_n8058;
  assign new_n8063 = n3852 & new_n8058;
  assign new_n8064 = n3851 & new_n8058;
  assign new_n8065 = n3850 & new_n8058;
  assign new_n8066 = n3849 & new_n8058;
  assign new_n8067 = new_n5524 & new_n8031;
  assign new_n8068 = ~new_n8067 & new_n8056;
  assign new_n8069 = n3848 & new_n8068;
  assign new_n8070 = n3847 & new_n8068;
  assign new_n8071 = n3846 & new_n8068;
  assign new_n8072 = n3845 & new_n8068;
  assign new_n8073 = n3844 & new_n8068;
  assign new_n8074 = n3843 & new_n8068;
  assign new_n8075 = n3842 & new_n8068;
  assign new_n8076 = n3841 & new_n8068;
  assign new_n8077 = new_n5485 & new_n6557;
  assign new_n8078 = new_n5434 & new_n8077;
  assign new_n8079 = new_n5430 & new_n8077;
  assign new_n8080 = ~new_n8078 & ~new_n8079;
  assign new_n8081 = new_n5438 & new_n8077;
  assign new_n8082 = ~new_n8081 & new_n8080;
  assign new_n8083 = n3904 & new_n8082;
  assign new_n8084 = n3903 & new_n8082;
  assign new_n8085 = n3902 & new_n8082;
  assign new_n8086 = n3901 & new_n8082;
  assign new_n8087 = n3900 & new_n8082;
  assign new_n8088 = n3899 & new_n8082;
  assign new_n8089 = n3898 & new_n8082;
  assign new_n8090 = n3897 & new_n8082;
  assign new_n8091 = new_n5500 & new_n8077;
  assign new_n8092 = ~new_n8091 & new_n8080;
  assign new_n8093 = n3896 & new_n8092;
  assign new_n8094 = n3895 & new_n8092;
  assign new_n8095 = n3894 & new_n8092;
  assign new_n8096 = n3893 & new_n8092;
  assign new_n8097 = n3892 & new_n8092;
  assign new_n8098 = n3891 & new_n8092;
  assign new_n8099 = n3890 & new_n8092;
  assign new_n8100 = n3889 & new_n8092;
  assign new_n8101 = new_n5433 & new_n8077;
  assign new_n8102 = ~new_n8079 & ~new_n8101;
  assign new_n8103 = new_n5513 & new_n8077;
  assign new_n8104 = ~new_n8103 & new_n8102;
  assign new_n8105 = n3888 & new_n8104;
  assign new_n8106 = n3887 & new_n8104;
  assign new_n8107 = n3886 & new_n8104;
  assign new_n8108 = n3885 & new_n8104;
  assign new_n8109 = n3884 & new_n8104;
  assign new_n8110 = n3883 & new_n8104;
  assign new_n8111 = n3882 & new_n8104;
  assign new_n8112 = n3881 & new_n8104;
  assign new_n8113 = new_n5524 & new_n8077;
  assign new_n8114 = ~new_n8113 & new_n8102;
  assign new_n8115 = n3880 & new_n8114;
  assign new_n8116 = n3879 & new_n8114;
  assign new_n8117 = n3878 & new_n8114;
  assign new_n8118 = n3877 & new_n8114;
  assign new_n8119 = n3876 & new_n8114;
  assign new_n8120 = n3875 & new_n8114;
  assign new_n8121 = n3874 & new_n8114;
  assign new_n8122 = n3873 & new_n8114;
  assign new_n8123 = new_n5537 & new_n6557;
  assign new_n8124 = new_n5434 & new_n8123;
  assign new_n8125 = new_n5430 & new_n8123;
  assign new_n8126 = ~new_n8124 & ~new_n8125;
  assign new_n8127 = new_n5438 & new_n8123;
  assign new_n8128 = ~new_n8127 & new_n8126;
  assign new_n8129 = n3936 & new_n8128;
  assign new_n8130 = n3935 & new_n8128;
  assign new_n8131 = n3934 & new_n8128;
  assign new_n8132 = n3933 & new_n8128;
  assign new_n8133 = n3932 & new_n8128;
  assign new_n8134 = n3931 & new_n8128;
  assign new_n8135 = n3930 & new_n8128;
  assign new_n8136 = n3929 & new_n8128;
  assign new_n8137 = new_n5500 & new_n8123;
  assign new_n8138 = ~new_n8137 & new_n8126;
  assign new_n8139 = n3928 & new_n8138;
  assign new_n8140 = n3927 & new_n8138;
  assign new_n8141 = n3926 & new_n8138;
  assign new_n8142 = n3925 & new_n8138;
  assign new_n8143 = n3924 & new_n8138;
  assign new_n8144 = n3923 & new_n8138;
  assign new_n8145 = n3922 & new_n8138;
  assign new_n8146 = n3921 & new_n8138;
  assign new_n8147 = new_n5433 & new_n8123;
  assign new_n8148 = ~new_n8125 & ~new_n8147;
  assign new_n8149 = new_n5513 & new_n8123;
  assign new_n8150 = ~new_n8149 & new_n8148;
  assign new_n8151 = n3920 & new_n8150;
  assign new_n8152 = n3919 & new_n8150;
  assign new_n8153 = n3918 & new_n8150;
  assign new_n8154 = n3917 & new_n8150;
  assign new_n8155 = n3916 & new_n8150;
  assign new_n8156 = n3915 & new_n8150;
  assign new_n8157 = n3914 & new_n8150;
  assign new_n8158 = n3913 & new_n8150;
  assign new_n8159 = new_n5524 & new_n8123;
  assign new_n8160 = ~new_n8159 & new_n8148;
  assign new_n8161 = n3912 & new_n8160;
  assign new_n8162 = n3911 & new_n8160;
  assign new_n8163 = n3910 & new_n8160;
  assign new_n8164 = n3909 & new_n8160;
  assign new_n8165 = n3908 & new_n8160;
  assign new_n8166 = n3907 & new_n8160;
  assign new_n8167 = n3906 & new_n8160;
  assign new_n8168 = n3905 & new_n8160;
  assign new_n8169 = new_n5245 & new_n6557;
  assign new_n8170 = new_n5434 & new_n8169;
  assign new_n8171 = new_n5430 & new_n8169;
  assign new_n8172 = ~new_n8170 & ~new_n8171;
  assign new_n8173 = new_n5438 & new_n8169;
  assign new_n8174 = ~new_n8173 & new_n8172;
  assign new_n8175 = n3968 & new_n8174;
  assign new_n8176 = n3967 & new_n8174;
  assign new_n8177 = n3966 & new_n8174;
  assign new_n8178 = n3965 & new_n8174;
  assign new_n8179 = n3964 & new_n8174;
  assign new_n8180 = n3963 & new_n8174;
  assign new_n8181 = n3962 & new_n8174;
  assign new_n8182 = n3961 & new_n8174;
  assign new_n8183 = new_n5500 & new_n8169;
  assign new_n8184 = ~new_n8183 & new_n8172;
  assign new_n8185 = n3960 & new_n8184;
  assign new_n8186 = n3959 & new_n8184;
  assign new_n8187 = n3958 & new_n8184;
  assign new_n8188 = n3957 & new_n8184;
  assign new_n8189 = n3956 & new_n8184;
  assign new_n8190 = n3955 & new_n8184;
  assign new_n8191 = n3954 & new_n8184;
  assign new_n8192 = n3953 & new_n8184;
  assign new_n8193 = new_n5433 & new_n8169;
  assign new_n8194 = ~new_n8171 & ~new_n8193;
  assign new_n8195 = new_n5513 & new_n8169;
  assign new_n8196 = ~new_n8195 & new_n8194;
  assign new_n8197 = n3952 & new_n8196;
  assign new_n8198 = n3951 & new_n8196;
  assign new_n8199 = n3950 & new_n8196;
  assign new_n8200 = n3949 & new_n8196;
  assign new_n8201 = n3948 & new_n8196;
  assign new_n8202 = n3947 & new_n8196;
  assign new_n8203 = n3946 & new_n8196;
  assign new_n8204 = n3945 & new_n8196;
  assign new_n8205 = new_n5524 & new_n8169;
  assign new_n8206 = ~new_n8205 & new_n8194;
  assign new_n8207 = n3944 & new_n8206;
  assign new_n8208 = n3943 & new_n8206;
  assign new_n8209 = n3942 & new_n8206;
  assign new_n8210 = n3941 & new_n8206;
  assign new_n8211 = n3940 & new_n8206;
  assign new_n8212 = n3939 & new_n8206;
  assign new_n8213 = n3938 & new_n8206;
  assign new_n8214 = n3937 & new_n8206;
  assign new_n8215 = new_n5423 & new_n6557;
  assign new_n8216 = new_n5434 & new_n8215;
  assign new_n8217 = new_n5430 & new_n8215;
  assign new_n8218 = ~new_n8216 & ~new_n8217;
  assign new_n8219 = new_n5438 & new_n8215;
  assign new_n8220 = ~new_n8219 & new_n8218;
  assign new_n8221 = n4000 & new_n8220;
  assign new_n8222 = n3999 & new_n8220;
  assign new_n8223 = n3998 & new_n8220;
  assign new_n8224 = n3997 & new_n8220;
  assign new_n8225 = n3996 & new_n8220;
  assign new_n8226 = n3995 & new_n8220;
  assign new_n8227 = n3994 & new_n8220;
  assign new_n8228 = n3993 & new_n8220;
  assign new_n8229 = new_n5500 & new_n8215;
  assign new_n8230 = ~new_n8229 & new_n8218;
  assign new_n8231 = n3992 & new_n8230;
  assign new_n8232 = n3991 & new_n8230;
  assign new_n8233 = n3990 & new_n8230;
  assign new_n8234 = n3989 & new_n8230;
  assign new_n8235 = n3988 & new_n8230;
  assign new_n8236 = n3987 & new_n8230;
  assign new_n8237 = n3986 & new_n8230;
  assign new_n8238 = n3985 & new_n8230;
  assign new_n8239 = new_n5433 & new_n8215;
  assign new_n8240 = ~new_n8217 & ~new_n8239;
  assign new_n8241 = new_n5513 & new_n8215;
  assign new_n8242 = ~new_n8241 & new_n8240;
  assign new_n8243 = n3984 & new_n8242;
  assign new_n8244 = n3983 & new_n8242;
  assign new_n8245 = n3982 & new_n8242;
  assign new_n8246 = n3981 & new_n8242;
  assign new_n8247 = n3980 & new_n8242;
  assign new_n8248 = n3979 & new_n8242;
  assign new_n8249 = n3978 & new_n8242;
  assign new_n8250 = n3977 & new_n8242;
  assign new_n8251 = new_n5524 & new_n8215;
  assign new_n8252 = ~new_n8251 & new_n8240;
  assign new_n8253 = n3976 & new_n8252;
  assign new_n8254 = n3975 & new_n8252;
  assign new_n8255 = n3974 & new_n8252;
  assign new_n8256 = n3973 & new_n8252;
  assign new_n8257 = n3972 & new_n8252;
  assign new_n8258 = n3971 & new_n8252;
  assign new_n8259 = n3970 & new_n8252;
  assign new_n8260 = n3969 & new_n8252;
  assign new_n8261 = new_n5484 & new_n6557;
  assign new_n8262 = new_n5434 & new_n8261;
  assign new_n8263 = new_n5430 & new_n8261;
  assign new_n8264 = ~new_n8262 & ~new_n8263;
  assign new_n8265 = new_n5438 & new_n8261;
  assign new_n8266 = ~new_n8265 & new_n8264;
  assign new_n8267 = n4032 & new_n8266;
  assign new_n8268 = n4031 & new_n8266;
  assign new_n8269 = n4030 & new_n8266;
  assign new_n8270 = n4029 & new_n8266;
  assign new_n8271 = n4028 & new_n8266;
  assign new_n8272 = n4027 & new_n8266;
  assign new_n8273 = n4026 & new_n8266;
  assign new_n8274 = n4025 & new_n8266;
  assign new_n8275 = new_n5500 & new_n8261;
  assign new_n8276 = ~new_n8275 & new_n8264;
  assign new_n8277 = n4024 & new_n8276;
  assign new_n8278 = n4023 & new_n8276;
  assign new_n8279 = n4022 & new_n8276;
  assign new_n8280 = n4021 & new_n8276;
  assign new_n8281 = n4020 & new_n8276;
  assign new_n8282 = n4019 & new_n8276;
  assign new_n8283 = n4018 & new_n8276;
  assign new_n8284 = n4017 & new_n8276;
  assign new_n8285 = new_n5433 & new_n8261;
  assign new_n8286 = ~new_n8263 & ~new_n8285;
  assign new_n8287 = new_n5513 & new_n8261;
  assign new_n8288 = ~new_n8287 & new_n8286;
  assign new_n8289 = n4016 & new_n8288;
  assign new_n8290 = n4015 & new_n8288;
  assign new_n8291 = n4014 & new_n8288;
  assign new_n8292 = n4013 & new_n8288;
  assign new_n8293 = n4012 & new_n8288;
  assign new_n8294 = n4011 & new_n8288;
  assign new_n8295 = n4010 & new_n8288;
  assign new_n8296 = n4009 & new_n8288;
  assign new_n8297 = new_n5524 & new_n8261;
  assign new_n8298 = ~new_n8297 & new_n8286;
  assign new_n8299 = n4008 & new_n8298;
  assign new_n8300 = n4007 & new_n8298;
  assign new_n8301 = n4006 & new_n8298;
  assign new_n8302 = n4005 & new_n8298;
  assign new_n8303 = n4004 & new_n8298;
  assign new_n8304 = n4003 & new_n8298;
  assign new_n8305 = n4002 & new_n8298;
  assign new_n8306 = n4001 & new_n8298;
  assign new_n8307 = new_n5536 & new_n6557;
  assign new_n8308 = new_n5434 & new_n8307;
  assign new_n8309 = new_n5430 & new_n8307;
  assign new_n8310 = ~new_n8308 & ~new_n8309;
  assign new_n8311 = new_n5438 & new_n8307;
  assign new_n8312 = ~new_n8311 & new_n8310;
  assign new_n8313 = n4064 & new_n8312;
  assign new_n8314 = n4063 & new_n8312;
  assign new_n8315 = n4062 & new_n8312;
  assign new_n8316 = n4061 & new_n8312;
  assign new_n8317 = n4060 & new_n8312;
  assign new_n8318 = n4059 & new_n8312;
  assign new_n8319 = n4058 & new_n8312;
  assign new_n8320 = n4057 & new_n8312;
  assign new_n8321 = new_n5500 & new_n8307;
  assign new_n8322 = ~new_n8321 & new_n8310;
  assign new_n8323 = n4056 & new_n8322;
  assign new_n8324 = n4055 & new_n8322;
  assign new_n8325 = n4054 & new_n8322;
  assign new_n8326 = n4053 & new_n8322;
  assign new_n8327 = n4052 & new_n8322;
  assign new_n8328 = n4051 & new_n8322;
  assign new_n8329 = n4050 & new_n8322;
  assign new_n8330 = n4049 & new_n8322;
  assign new_n8331 = new_n5433 & new_n8307;
  assign new_n8332 = ~new_n8309 & ~new_n8331;
  assign new_n8333 = new_n5513 & new_n8307;
  assign new_n8334 = ~new_n8333 & new_n8332;
  assign new_n8335 = n4048 & new_n8334;
  assign new_n8336 = n4047 & new_n8334;
  assign new_n8337 = n4046 & new_n8334;
  assign new_n8338 = n4045 & new_n8334;
  assign new_n8339 = n4044 & new_n8334;
  assign new_n8340 = n4043 & new_n8334;
  assign new_n8341 = n4042 & new_n8334;
  assign new_n8342 = n4041 & new_n8334;
  assign new_n8343 = new_n5524 & new_n8307;
  assign new_n8344 = ~new_n8343 & new_n8332;
  assign new_n8345 = n4040 & new_n8344;
  assign new_n8346 = n4039 & new_n8344;
  assign new_n8347 = n4038 & new_n8344;
  assign new_n8348 = n4037 & new_n8344;
  assign new_n8349 = n4036 & new_n8344;
  assign new_n8350 = n4035 & new_n8344;
  assign new_n8351 = n4034 & new_n8344;
  assign new_n8352 = n4033 & new_n8344;
  assign new_n8353 = new_n5246 & new_n6557;
  assign new_n8354 = new_n5430 & new_n8353;
  assign new_n8355 = new_n5434 & new_n8353;
  assign new_n8356 = ~new_n8354 & ~new_n8355;
  assign new_n8357 = new_n5438 & new_n8353;
  assign new_n8358 = ~new_n8357 & new_n8356;
  assign new_n8359 = n4096 & new_n8358;
  assign new_n8360 = n4095 & new_n8358;
  assign new_n8361 = n4094 & new_n8358;
  assign new_n8362 = n4093 & new_n8358;
  assign new_n8363 = n4092 & new_n8358;
  assign new_n8364 = n4091 & new_n8358;
  assign new_n8365 = n4090 & new_n8358;
  assign new_n8366 = n4089 & new_n8358;
  assign new_n8367 = new_n5500 & new_n8353;
  assign new_n8368 = ~new_n8367 & new_n8356;
  assign new_n8369 = n4088 & new_n8368;
  assign new_n8370 = n4087 & new_n8368;
  assign new_n8371 = n4086 & new_n8368;
  assign new_n8372 = n4085 & new_n8368;
  assign new_n8373 = n4084 & new_n8368;
  assign new_n8374 = n4083 & new_n8368;
  assign new_n8375 = n4082 & new_n8368;
  assign new_n8376 = n4081 & new_n8368;
  assign new_n8377 = new_n5433 & new_n8353;
  assign new_n8378 = ~new_n8354 & ~new_n8377;
  assign new_n8379 = new_n5513 & new_n8353;
  assign new_n8380 = ~new_n8379 & new_n8378;
  assign new_n8381 = n4080 & new_n8380;
  assign new_n8382 = n4079 & new_n8380;
  assign new_n8383 = n4078 & new_n8380;
  assign new_n8384 = n4077 & new_n8380;
  assign new_n8385 = n4076 & new_n8380;
  assign new_n8386 = n4075 & new_n8380;
  assign new_n8387 = n4074 & new_n8380;
  assign new_n8388 = n4073 & new_n8380;
  assign new_n8389 = new_n5524 & new_n8353;
  assign new_n8390 = ~new_n8389 & new_n8378;
  assign new_n8391 = n4072 & new_n8390;
  assign new_n8392 = n4071 & new_n8390;
  assign new_n8393 = n4070 & new_n8390;
  assign new_n8394 = n4069 & new_n8390;
  assign new_n8395 = n4068 & new_n8390;
  assign new_n8396 = n4067 & new_n8390;
  assign new_n8397 = n4066 & new_n8390;
  assign new_n8398 = n4065 & new_n8390;
  assign new_n8399 = new_n5429 ^ new_n4151;
  assign new_n8400 = ~new_n8399 & n2029;
  assign new_n8401 = ~n2025 & ~n2029;
  assign new_n8402 = ~new_n8401 & new_n4266;
  assign new_n8403 = ~n2034 & n2025;
  assign new_n8404 = ~new_n8403 & new_n8402;
  assign new_n8405 = ~new_n8400 & ~new_n8404;
  assign new_n8406 = n2034 & new_n4114;
  assign new_n8407 = new_n4112 ^ n2047;
  assign new_n8408 = ~new_n8406 & new_n8407;
  assign new_n8409 = ~new_n8408 & new_n4269;
  assign new_n8410 = ~new_n4293 & n2034;
  assign new_n8411 = ~new_n4271 & new_n8410;
  assign new_n8412 = ~new_n8409 & ~new_n8411;
  assign new_n8413 = ~new_n4276 & new_n4110;
  assign new_n8414 = ~new_n4109 & ~new_n8413;
  assign new_n8415 = ~n2043 & ~n2045;
  assign new_n8416 = ~new_n4273 & new_n8415;
  assign new_n8417 = ~new_n8416 & new_n8414;
  assign new_n8418 = ~new_n8417 & n2034;
  assign new_n8419 = ~new_n8418 & new_n8412;
  assign new_n8420 = ~new_n4107 & ~new_n8419;
  assign new_n8421 = n2028 & new_n4286;
  assign new_n8422 = new_n8421 ^ new_n4136;
  assign new_n8423 = ~new_n8420 & ~new_n8422;
  assign new_n8424 = ~new_n8423 & new_n4118;
  assign new_n8425 = ~new_n4132 & n2029;
  assign new_n8426 = ~new_n8424 & ~new_n8425;
  assign new_n8427 = new_n8405 & new_n8426;
  assign new_n8428 = ~new_n8399 & n2028;
  assign new_n8429 = ~n2025 & ~n2028;
  assign new_n8430 = ~new_n8429 & new_n4266;
  assign new_n8431 = ~n2033 & n2025;
  assign new_n8432 = ~new_n8431 & new_n8430;
  assign new_n8433 = ~new_n8428 & ~new_n8432;
  assign new_n8434 = n2033 & new_n4269;
  assign new_n8435 = new_n4114 & new_n8434;
  assign new_n8436 = ~new_n4293 & n2033;
  assign new_n8437 = ~new_n4271 & new_n8436;
  assign new_n8438 = ~new_n8435 & ~new_n8437;
  assign new_n8439 = ~new_n8417 & n2033;
  assign new_n8440 = ~new_n8439 & new_n8438;
  assign new_n8441 = ~new_n4107 & ~new_n8440;
  assign new_n8442 = ~new_n8422 & ~new_n8441;
  assign new_n8443 = ~new_n8442 & new_n4118;
  assign new_n8444 = ~new_n4132 & n2028;
  assign new_n8445 = ~new_n8443 & ~new_n8444;
  assign new_n8446 = new_n8433 & new_n8445;
  assign new_n8447 = ~new_n8427 & ~new_n8446;
  assign new_n8448 = new_n8447 ^ new_n8446;
  assign new_n8449 = new_n8448 ^ new_n8427;
  assign new_n8450 = ~new_n8399 & n2032;
  assign new_n8451 = ~n2025 & ~n2032;
  assign new_n8452 = ~new_n8451 & new_n4266;
  assign new_n8453 = ~n2037 & n2025;
  assign new_n8454 = ~new_n8453 & new_n8452;
  assign new_n8455 = ~new_n8450 & ~new_n8454;
  assign new_n8456 = n2037 & new_n4269;
  assign new_n8457 = new_n4114 & new_n8456;
  assign new_n8458 = ~new_n4293 & n2037;
  assign new_n8459 = ~new_n4271 & new_n8458;
  assign new_n8460 = ~new_n8457 & ~new_n8459;
  assign new_n8461 = ~new_n8417 & n2037;
  assign new_n8462 = ~new_n8461 & new_n8460;
  assign new_n8463 = ~new_n4107 & ~new_n8462;
  assign new_n8464 = ~new_n8422 & ~new_n8463;
  assign new_n8465 = ~new_n8464 & new_n4118;
  assign new_n8466 = ~new_n4132 & n2032;
  assign new_n8467 = ~new_n8465 & ~new_n8466;
  assign new_n8468 = new_n8455 & new_n8467;
  assign new_n8469 = ~new_n8399 & n2031;
  assign new_n8470 = ~n2025 & ~n2031;
  assign new_n8471 = ~new_n8470 & new_n4266;
  assign new_n8472 = ~n2036 & n2025;
  assign new_n8473 = ~new_n8472 & new_n8471;
  assign new_n8474 = ~new_n8469 & ~new_n8473;
  assign new_n8475 = n2036 & new_n4114;
  assign new_n8476 = ~new_n8475 & new_n8407;
  assign new_n8477 = ~new_n8476 & new_n4269;
  assign new_n8478 = ~new_n4293 & n2036;
  assign new_n8479 = ~new_n4271 & new_n8478;
  assign new_n8480 = ~new_n8477 & ~new_n8479;
  assign new_n8481 = ~new_n8417 & n2036;
  assign new_n8482 = ~new_n8481 & new_n8480;
  assign new_n8483 = ~new_n4107 & ~new_n8482;
  assign new_n8484 = ~new_n8422 & ~new_n8483;
  assign new_n8485 = ~new_n8484 & new_n4118;
  assign new_n8486 = ~new_n4132 & n2031;
  assign new_n8487 = ~new_n8485 & ~new_n8486;
  assign new_n8488 = new_n8474 & new_n8487;
  assign new_n8489 = new_n8468 & new_n8488;
  assign new_n8490 = new_n8489 ^ new_n8468;
  assign new_n8491 = new_n8490 ^ new_n8488;
  assign new_n8492 = new_n8491 ^ new_n8468;
  assign new_n8493 = ~new_n8399 & n2030;
  assign new_n8494 = ~n2025 & ~n2030;
  assign new_n8495 = ~new_n8494 & new_n4266;
  assign new_n8496 = ~n2035 & n2025;
  assign new_n8497 = ~new_n8496 & new_n8495;
  assign new_n8498 = ~new_n8493 & ~new_n8497;
  assign new_n8499 = n2035 & new_n4114;
  assign new_n8500 = ~new_n8499 & new_n8407;
  assign new_n8501 = ~new_n8500 & new_n4269;
  assign new_n8502 = ~new_n4293 & n2035;
  assign new_n8503 = ~new_n4271 & new_n8502;
  assign new_n8504 = ~new_n8501 & ~new_n8503;
  assign new_n8505 = ~new_n8417 & n2035;
  assign new_n8506 = ~new_n8505 & new_n8504;
  assign new_n8507 = ~new_n4107 & ~new_n8506;
  assign new_n8508 = ~new_n8422 & ~new_n8507;
  assign new_n8509 = ~new_n8508 & new_n4118;
  assign new_n8510 = ~new_n4132 & n2030;
  assign new_n8511 = ~new_n8509 & ~new_n8510;
  assign new_n8512 = new_n8498 & new_n8511;
  assign new_n8513 = ~new_n8512 & new_n8492;
  assign new_n8514 = new_n8513 ^ new_n8492;
  assign new_n8515 = ~new_n8449 & new_n8514;
  assign new_n8516 = ~new_n5207 & n2080;
  assign new_n8517 = n2112 & new_n5207;
  assign new_n8518 = ~new_n8516 & ~new_n8517;
  assign new_n8519 = ~new_n5243 & ~new_n8518;
  assign new_n8520 = ~new_n5207 & n2144;
  assign new_n8521 = n2176 & new_n5207;
  assign new_n8522 = ~new_n8520 & ~new_n8521;
  assign new_n8523 = ~new_n8522 & new_n5243;
  assign new_n8524 = ~new_n8519 & ~new_n8523;
  assign new_n8525 = ~new_n5170 & ~new_n8524;
  assign new_n8526 = ~new_n5207 & n2208;
  assign new_n8527 = n2240 & new_n5207;
  assign new_n8528 = ~new_n8526 & ~new_n8527;
  assign new_n8529 = ~new_n5243 & ~new_n8528;
  assign new_n8530 = ~new_n5207 & n2272;
  assign new_n8531 = n2304 & new_n5207;
  assign new_n8532 = ~new_n8530 & ~new_n8531;
  assign new_n8533 = ~new_n8532 & new_n5243;
  assign new_n8534 = ~new_n8529 & ~new_n8533;
  assign new_n8535 = ~new_n8534 & new_n5170;
  assign new_n8536 = ~new_n8525 & ~new_n8535;
  assign new_n8537 = ~new_n5139 & ~new_n8536;
  assign new_n8538 = ~new_n5207 & n2336;
  assign new_n8539 = n2368 & new_n5207;
  assign new_n8540 = ~new_n8538 & ~new_n8539;
  assign new_n8541 = ~new_n5243 & ~new_n8540;
  assign new_n8542 = ~new_n5207 & n2400;
  assign new_n8543 = n2432 & new_n5207;
  assign new_n8544 = ~new_n8542 & ~new_n8543;
  assign new_n8545 = ~new_n8544 & new_n5243;
  assign new_n8546 = ~new_n8541 & ~new_n8545;
  assign new_n8547 = ~new_n5170 & ~new_n8546;
  assign new_n8548 = ~new_n5207 & n2464;
  assign new_n8549 = n2496 & new_n5207;
  assign new_n8550 = ~new_n8548 & ~new_n8549;
  assign new_n8551 = ~new_n5243 & ~new_n8550;
  assign new_n8552 = ~new_n5207 & n2528;
  assign new_n8553 = n2560 & new_n5207;
  assign new_n8554 = ~new_n8552 & ~new_n8553;
  assign new_n8555 = ~new_n8554 & new_n5243;
  assign new_n8556 = ~new_n8551 & ~new_n8555;
  assign new_n8557 = ~new_n8556 & new_n5170;
  assign new_n8558 = ~new_n8547 & ~new_n8557;
  assign new_n8559 = ~new_n8558 & new_n5139;
  assign new_n8560 = ~new_n8537 & ~new_n8559;
  assign new_n8561 = ~new_n5011 & ~new_n8560;
  assign new_n8562 = ~new_n5207 & n2592;
  assign new_n8563 = n2624 & new_n5207;
  assign new_n8564 = ~new_n8562 & ~new_n8563;
  assign new_n8565 = ~new_n5243 & ~new_n8564;
  assign new_n8566 = ~new_n5207 & n2656;
  assign new_n8567 = n2688 & new_n5207;
  assign new_n8568 = ~new_n8566 & ~new_n8567;
  assign new_n8569 = ~new_n8568 & new_n5243;
  assign new_n8570 = ~new_n8565 & ~new_n8569;
  assign new_n8571 = ~new_n5170 & ~new_n8570;
  assign new_n8572 = ~new_n5207 & n2720;
  assign new_n8573 = n2752 & new_n5207;
  assign new_n8574 = ~new_n8572 & ~new_n8573;
  assign new_n8575 = ~new_n5243 & ~new_n8574;
  assign new_n8576 = ~new_n5207 & n2784;
  assign new_n8577 = n2816 & new_n5207;
  assign new_n8578 = ~new_n8576 & ~new_n8577;
  assign new_n8579 = ~new_n8578 & new_n5243;
  assign new_n8580 = ~new_n8575 & ~new_n8579;
  assign new_n8581 = ~new_n8580 & new_n5170;
  assign new_n8582 = ~new_n8571 & ~new_n8581;
  assign new_n8583 = ~new_n5139 & ~new_n8582;
  assign new_n8584 = ~new_n5207 & n2848;
  assign new_n8585 = n2880 & new_n5207;
  assign new_n8586 = ~new_n8584 & ~new_n8585;
  assign new_n8587 = ~new_n5243 & ~new_n8586;
  assign new_n8588 = ~new_n5207 & n2912;
  assign new_n8589 = n2944 & new_n5207;
  assign new_n8590 = ~new_n8588 & ~new_n8589;
  assign new_n8591 = ~new_n8590 & new_n5243;
  assign new_n8592 = ~new_n8587 & ~new_n8591;
  assign new_n8593 = ~new_n5170 & ~new_n8592;
  assign new_n8594 = ~new_n5207 & n2976;
  assign new_n8595 = n3008 & new_n5207;
  assign new_n8596 = ~new_n8594 & ~new_n8595;
  assign new_n8597 = ~new_n5243 & ~new_n8596;
  assign new_n8598 = ~new_n5207 & n3040;
  assign new_n8599 = n3072 & new_n5207;
  assign new_n8600 = ~new_n8598 & ~new_n8599;
  assign new_n8601 = ~new_n8600 & new_n5243;
  assign new_n8602 = ~new_n8597 & ~new_n8601;
  assign new_n8603 = ~new_n8602 & new_n5170;
  assign new_n8604 = ~new_n8593 & ~new_n8603;
  assign new_n8605 = ~new_n8604 & new_n5139;
  assign new_n8606 = ~new_n8583 & ~new_n8605;
  assign new_n8607 = ~new_n8606 & new_n5011;
  assign new_n8608 = ~new_n8561 & ~new_n8607;
  assign new_n8609 = ~new_n5031 & ~new_n8608;
  assign new_n8610 = ~new_n5207 & n3104;
  assign new_n8611 = n3136 & new_n5207;
  assign new_n8612 = ~new_n8610 & ~new_n8611;
  assign new_n8613 = ~new_n5243 & ~new_n8612;
  assign new_n8614 = ~new_n5207 & n3168;
  assign new_n8615 = n3200 & new_n5207;
  assign new_n8616 = ~new_n8614 & ~new_n8615;
  assign new_n8617 = ~new_n8616 & new_n5243;
  assign new_n8618 = ~new_n8613 & ~new_n8617;
  assign new_n8619 = ~new_n5170 & ~new_n8618;
  assign new_n8620 = ~new_n5207 & n3232;
  assign new_n8621 = n3264 & new_n5207;
  assign new_n8622 = ~new_n8620 & ~new_n8621;
  assign new_n8623 = ~new_n5243 & ~new_n8622;
  assign new_n8624 = ~new_n5207 & n3296;
  assign new_n8625 = n3328 & new_n5207;
  assign new_n8626 = ~new_n8624 & ~new_n8625;
  assign new_n8627 = ~new_n8626 & new_n5243;
  assign new_n8628 = ~new_n8623 & ~new_n8627;
  assign new_n8629 = ~new_n8628 & new_n5170;
  assign new_n8630 = ~new_n8619 & ~new_n8629;
  assign new_n8631 = ~new_n5139 & ~new_n8630;
  assign new_n8632 = ~new_n5207 & n3360;
  assign new_n8633 = n3392 & new_n5207;
  assign new_n8634 = ~new_n8632 & ~new_n8633;
  assign new_n8635 = ~new_n5243 & ~new_n8634;
  assign new_n8636 = ~new_n5207 & n3424;
  assign new_n8637 = n3456 & new_n5207;
  assign new_n8638 = ~new_n8636 & ~new_n8637;
  assign new_n8639 = ~new_n8638 & new_n5243;
  assign new_n8640 = ~new_n8635 & ~new_n8639;
  assign new_n8641 = ~new_n5170 & ~new_n8640;
  assign new_n8642 = ~new_n5207 & n3488;
  assign new_n8643 = n3520 & new_n5207;
  assign new_n8644 = ~new_n8642 & ~new_n8643;
  assign new_n8645 = ~new_n5243 & ~new_n8644;
  assign new_n8646 = ~new_n5207 & n3552;
  assign new_n8647 = n3584 & new_n5207;
  assign new_n8648 = ~new_n8646 & ~new_n8647;
  assign new_n8649 = ~new_n8648 & new_n5243;
  assign new_n8650 = ~new_n8645 & ~new_n8649;
  assign new_n8651 = ~new_n8650 & new_n5170;
  assign new_n8652 = ~new_n8641 & ~new_n8651;
  assign new_n8653 = ~new_n8652 & new_n5139;
  assign new_n8654 = ~new_n8631 & ~new_n8653;
  assign new_n8655 = ~new_n5011 & ~new_n8654;
  assign new_n8656 = ~new_n5207 & n3616;
  assign new_n8657 = n3648 & new_n5207;
  assign new_n8658 = ~new_n8656 & ~new_n8657;
  assign new_n8659 = ~new_n5243 & ~new_n8658;
  assign new_n8660 = ~new_n5207 & n3680;
  assign new_n8661 = n3712 & new_n5207;
  assign new_n8662 = ~new_n8660 & ~new_n8661;
  assign new_n8663 = ~new_n8662 & new_n5243;
  assign new_n8664 = ~new_n8659 & ~new_n8663;
  assign new_n8665 = ~new_n5170 & ~new_n8664;
  assign new_n8666 = ~new_n5207 & n3744;
  assign new_n8667 = n3776 & new_n5207;
  assign new_n8668 = ~new_n8666 & ~new_n8667;
  assign new_n8669 = ~new_n5243 & ~new_n8668;
  assign new_n8670 = ~new_n5207 & n3808;
  assign new_n8671 = n3840 & new_n5207;
  assign new_n8672 = ~new_n8670 & ~new_n8671;
  assign new_n8673 = ~new_n8672 & new_n5243;
  assign new_n8674 = ~new_n8669 & ~new_n8673;
  assign new_n8675 = ~new_n8674 & new_n5170;
  assign new_n8676 = ~new_n8665 & ~new_n8675;
  assign new_n8677 = ~new_n5139 & ~new_n8676;
  assign new_n8678 = ~new_n5207 & n3872;
  assign new_n8679 = n3904 & new_n5207;
  assign new_n8680 = ~new_n8678 & ~new_n8679;
  assign new_n8681 = ~new_n5243 & ~new_n8680;
  assign new_n8682 = ~new_n5207 & n3936;
  assign new_n8683 = n3968 & new_n5207;
  assign new_n8684 = ~new_n8682 & ~new_n8683;
  assign new_n8685 = ~new_n8684 & new_n5243;
  assign new_n8686 = ~new_n8681 & ~new_n8685;
  assign new_n8687 = ~new_n5170 & ~new_n8686;
  assign new_n8688 = ~new_n5207 & n4000;
  assign new_n8689 = n4032 & new_n5207;
  assign new_n8690 = ~new_n8688 & ~new_n8689;
  assign new_n8691 = ~new_n5243 & ~new_n8690;
  assign new_n8692 = ~new_n5207 & n4064;
  assign new_n8693 = n4096 & new_n5207;
  assign new_n8694 = ~new_n8692 & ~new_n8693;
  assign new_n8695 = ~new_n8694 & new_n5243;
  assign new_n8696 = ~new_n8691 & ~new_n8695;
  assign new_n8697 = ~new_n8696 & new_n5170;
  assign new_n8698 = ~new_n8687 & ~new_n8697;
  assign new_n8699 = ~new_n8698 & new_n5139;
  assign new_n8700 = ~new_n8677 & ~new_n8699;
  assign new_n8701 = ~new_n8700 & new_n5011;
  assign new_n8702 = ~new_n8655 & ~new_n8701;
  assign new_n8703 = ~new_n8702 & new_n5031;
  assign new_n8704 = ~new_n8609 & ~new_n8703;
  assign new_n8705 = ~new_n8704 & new_n5077;
  assign new_n8706 = ~new_n5207 & n2064;
  assign new_n8707 = n2096 & new_n5207;
  assign new_n8708 = ~new_n8706 & ~new_n8707;
  assign new_n8709 = ~new_n5243 & ~new_n8708;
  assign new_n8710 = ~new_n5207 & n2128;
  assign new_n8711 = n2160 & new_n5207;
  assign new_n8712 = ~new_n8710 & ~new_n8711;
  assign new_n8713 = ~new_n8712 & new_n5243;
  assign new_n8714 = ~new_n8709 & ~new_n8713;
  assign new_n8715 = ~new_n5170 & ~new_n8714;
  assign new_n8716 = ~new_n5207 & n2192;
  assign new_n8717 = n2224 & new_n5207;
  assign new_n8718 = ~new_n8716 & ~new_n8717;
  assign new_n8719 = ~new_n5243 & ~new_n8718;
  assign new_n8720 = ~new_n5207 & n2256;
  assign new_n8721 = n2288 & new_n5207;
  assign new_n8722 = ~new_n8720 & ~new_n8721;
  assign new_n8723 = ~new_n8722 & new_n5243;
  assign new_n8724 = ~new_n8719 & ~new_n8723;
  assign new_n8725 = ~new_n8724 & new_n5170;
  assign new_n8726 = ~new_n8715 & ~new_n8725;
  assign new_n8727 = ~new_n5139 & ~new_n8726;
  assign new_n8728 = ~new_n5207 & n2320;
  assign new_n8729 = n2352 & new_n5207;
  assign new_n8730 = ~new_n8728 & ~new_n8729;
  assign new_n8731 = ~new_n5243 & ~new_n8730;
  assign new_n8732 = ~new_n5207 & n2384;
  assign new_n8733 = n2416 & new_n5207;
  assign new_n8734 = ~new_n8732 & ~new_n8733;
  assign new_n8735 = ~new_n8734 & new_n5243;
  assign new_n8736 = ~new_n8731 & ~new_n8735;
  assign new_n8737 = ~new_n5170 & ~new_n8736;
  assign new_n8738 = ~new_n5207 & n2448;
  assign new_n8739 = n2480 & new_n5207;
  assign new_n8740 = ~new_n8738 & ~new_n8739;
  assign new_n8741 = ~new_n5243 & ~new_n8740;
  assign new_n8742 = ~new_n5207 & n2512;
  assign new_n8743 = n2544 & new_n5207;
  assign new_n8744 = ~new_n8742 & ~new_n8743;
  assign new_n8745 = ~new_n8744 & new_n5243;
  assign new_n8746 = ~new_n8741 & ~new_n8745;
  assign new_n8747 = ~new_n8746 & new_n5170;
  assign new_n8748 = ~new_n8737 & ~new_n8747;
  assign new_n8749 = ~new_n8748 & new_n5139;
  assign new_n8750 = ~new_n8727 & ~new_n8749;
  assign new_n8751 = ~new_n5011 & ~new_n8750;
  assign new_n8752 = ~new_n5207 & n2576;
  assign new_n8753 = n2608 & new_n5207;
  assign new_n8754 = ~new_n8752 & ~new_n8753;
  assign new_n8755 = ~new_n5243 & ~new_n8754;
  assign new_n8756 = ~new_n5207 & n2640;
  assign new_n8757 = n2672 & new_n5207;
  assign new_n8758 = ~new_n8756 & ~new_n8757;
  assign new_n8759 = ~new_n8758 & new_n5243;
  assign new_n8760 = ~new_n8755 & ~new_n8759;
  assign new_n8761 = ~new_n5170 & ~new_n8760;
  assign new_n8762 = ~new_n5207 & n2704;
  assign new_n8763 = n2736 & new_n5207;
  assign new_n8764 = ~new_n8762 & ~new_n8763;
  assign new_n8765 = ~new_n5243 & ~new_n8764;
  assign new_n8766 = ~new_n5207 & n2768;
  assign new_n8767 = n2800 & new_n5207;
  assign new_n8768 = ~new_n8766 & ~new_n8767;
  assign new_n8769 = ~new_n8768 & new_n5243;
  assign new_n8770 = ~new_n8765 & ~new_n8769;
  assign new_n8771 = ~new_n8770 & new_n5170;
  assign new_n8772 = ~new_n8761 & ~new_n8771;
  assign new_n8773 = ~new_n5139 & ~new_n8772;
  assign new_n8774 = ~new_n5207 & n2832;
  assign new_n8775 = n2864 & new_n5207;
  assign new_n8776 = ~new_n8774 & ~new_n8775;
  assign new_n8777 = ~new_n5243 & ~new_n8776;
  assign new_n8778 = ~new_n5207 & n2896;
  assign new_n8779 = n2928 & new_n5207;
  assign new_n8780 = ~new_n8778 & ~new_n8779;
  assign new_n8781 = ~new_n8780 & new_n5243;
  assign new_n8782 = ~new_n8777 & ~new_n8781;
  assign new_n8783 = ~new_n5170 & ~new_n8782;
  assign new_n8784 = ~new_n5207 & n2960;
  assign new_n8785 = n2992 & new_n5207;
  assign new_n8786 = ~new_n8784 & ~new_n8785;
  assign new_n8787 = ~new_n5243 & ~new_n8786;
  assign new_n8788 = ~new_n5207 & n3024;
  assign new_n8789 = n3056 & new_n5207;
  assign new_n8790 = ~new_n8788 & ~new_n8789;
  assign new_n8791 = ~new_n8790 & new_n5243;
  assign new_n8792 = ~new_n8787 & ~new_n8791;
  assign new_n8793 = ~new_n8792 & new_n5170;
  assign new_n8794 = ~new_n8783 & ~new_n8793;
  assign new_n8795 = ~new_n8794 & new_n5139;
  assign new_n8796 = ~new_n8773 & ~new_n8795;
  assign new_n8797 = ~new_n8796 & new_n5011;
  assign new_n8798 = ~new_n8751 & ~new_n8797;
  assign new_n8799 = ~new_n5031 & ~new_n8798;
  assign new_n8800 = ~new_n5207 & n3088;
  assign new_n8801 = n3120 & new_n5207;
  assign new_n8802 = ~new_n8800 & ~new_n8801;
  assign new_n8803 = ~new_n5243 & ~new_n8802;
  assign new_n8804 = ~new_n5207 & n3152;
  assign new_n8805 = n3184 & new_n5207;
  assign new_n8806 = ~new_n8804 & ~new_n8805;
  assign new_n8807 = ~new_n8806 & new_n5243;
  assign new_n8808 = ~new_n8803 & ~new_n8807;
  assign new_n8809 = ~new_n5170 & ~new_n8808;
  assign new_n8810 = ~new_n5207 & n3216;
  assign new_n8811 = n3248 & new_n5207;
  assign new_n8812 = ~new_n8810 & ~new_n8811;
  assign new_n8813 = ~new_n5243 & ~new_n8812;
  assign new_n8814 = ~new_n5207 & n3280;
  assign new_n8815 = n3312 & new_n5207;
  assign new_n8816 = ~new_n8814 & ~new_n8815;
  assign new_n8817 = ~new_n8816 & new_n5243;
  assign new_n8818 = ~new_n8813 & ~new_n8817;
  assign new_n8819 = ~new_n8818 & new_n5170;
  assign new_n8820 = ~new_n8809 & ~new_n8819;
  assign new_n8821 = ~new_n5139 & ~new_n8820;
  assign new_n8822 = ~new_n5207 & n3344;
  assign new_n8823 = n3376 & new_n5207;
  assign new_n8824 = ~new_n8822 & ~new_n8823;
  assign new_n8825 = ~new_n5243 & ~new_n8824;
  assign new_n8826 = ~new_n5207 & n3408;
  assign new_n8827 = n3440 & new_n5207;
  assign new_n8828 = ~new_n8826 & ~new_n8827;
  assign new_n8829 = ~new_n8828 & new_n5243;
  assign new_n8830 = ~new_n8825 & ~new_n8829;
  assign new_n8831 = ~new_n5170 & ~new_n8830;
  assign new_n8832 = ~new_n5207 & n3472;
  assign new_n8833 = n3504 & new_n5207;
  assign new_n8834 = ~new_n8832 & ~new_n8833;
  assign new_n8835 = ~new_n5243 & ~new_n8834;
  assign new_n8836 = ~new_n5207 & n3536;
  assign new_n8837 = n3568 & new_n5207;
  assign new_n8838 = ~new_n8836 & ~new_n8837;
  assign new_n8839 = ~new_n8838 & new_n5243;
  assign new_n8840 = ~new_n8835 & ~new_n8839;
  assign new_n8841 = ~new_n8840 & new_n5170;
  assign new_n8842 = ~new_n8831 & ~new_n8841;
  assign new_n8843 = ~new_n8842 & new_n5139;
  assign new_n8844 = ~new_n8821 & ~new_n8843;
  assign new_n8845 = ~new_n5011 & ~new_n8844;
  assign new_n8846 = ~new_n5207 & n3600;
  assign new_n8847 = n3632 & new_n5207;
  assign new_n8848 = ~new_n8846 & ~new_n8847;
  assign new_n8849 = ~new_n5243 & ~new_n8848;
  assign new_n8850 = ~new_n5207 & n3664;
  assign new_n8851 = n3696 & new_n5207;
  assign new_n8852 = ~new_n8850 & ~new_n8851;
  assign new_n8853 = ~new_n8852 & new_n5243;
  assign new_n8854 = ~new_n8849 & ~new_n8853;
  assign new_n8855 = ~new_n5170 & ~new_n8854;
  assign new_n8856 = ~new_n5207 & n3728;
  assign new_n8857 = n3760 & new_n5207;
  assign new_n8858 = ~new_n8856 & ~new_n8857;
  assign new_n8859 = ~new_n5243 & ~new_n8858;
  assign new_n8860 = ~new_n5207 & n3792;
  assign new_n8861 = n3824 & new_n5207;
  assign new_n8862 = ~new_n8860 & ~new_n8861;
  assign new_n8863 = ~new_n8862 & new_n5243;
  assign new_n8864 = ~new_n8859 & ~new_n8863;
  assign new_n8865 = ~new_n8864 & new_n5170;
  assign new_n8866 = ~new_n8855 & ~new_n8865;
  assign new_n8867 = ~new_n5139 & ~new_n8866;
  assign new_n8868 = ~new_n5207 & n3856;
  assign new_n8869 = n3888 & new_n5207;
  assign new_n8870 = ~new_n8868 & ~new_n8869;
  assign new_n8871 = ~new_n5243 & ~new_n8870;
  assign new_n8872 = ~new_n5207 & n3920;
  assign new_n8873 = n3952 & new_n5207;
  assign new_n8874 = ~new_n8872 & ~new_n8873;
  assign new_n8875 = ~new_n8874 & new_n5243;
  assign new_n8876 = ~new_n8871 & ~new_n8875;
  assign new_n8877 = ~new_n5170 & ~new_n8876;
  assign new_n8878 = ~new_n5207 & n3984;
  assign new_n8879 = n4016 & new_n5207;
  assign new_n8880 = ~new_n8878 & ~new_n8879;
  assign new_n8881 = ~new_n5243 & ~new_n8880;
  assign new_n8882 = ~new_n5207 & n4048;
  assign new_n8883 = n4080 & new_n5207;
  assign new_n8884 = ~new_n8882 & ~new_n8883;
  assign new_n8885 = ~new_n8884 & new_n5243;
  assign new_n8886 = ~new_n8881 & ~new_n8885;
  assign new_n8887 = ~new_n8886 & new_n5170;
  assign new_n8888 = ~new_n8877 & ~new_n8887;
  assign new_n8889 = ~new_n8888 & new_n5139;
  assign new_n8890 = ~new_n8867 & ~new_n8889;
  assign new_n8891 = ~new_n8890 & new_n5011;
  assign new_n8892 = ~new_n8845 & ~new_n8891;
  assign new_n8893 = ~new_n8892 & new_n5031;
  assign new_n8894 = ~new_n8799 & ~new_n8893;
  assign new_n8895 = ~new_n5077 & ~new_n8894;
  assign new_n8896 = ~new_n8705 & ~new_n8895;
  assign new_n8897 = ~new_n4099 & new_n4142;
  assign new_n8898 = new_n4151 ^ new_n4149;
  assign new_n8899 = new_n8898 ^ new_n4144;
  assign new_n8900 = ~new_n8899 & new_n8897;
  assign new_n8901 = new_n8900 ^ new_n8897;
  assign new_n8902 = new_n8901 ^ new_n8898;
  assign new_n8903 = ~new_n8896 & new_n8902;
  assign new_n8904 = ~new_n5207 & n2056;
  assign new_n8905 = n2088 & new_n5207;
  assign new_n8906 = ~new_n8904 & ~new_n8905;
  assign new_n8907 = ~new_n5243 & ~new_n8906;
  assign new_n8908 = ~new_n5207 & n2120;
  assign new_n8909 = n2152 & new_n5207;
  assign new_n8910 = ~new_n8908 & ~new_n8909;
  assign new_n8911 = ~new_n8910 & new_n5243;
  assign new_n8912 = ~new_n8907 & ~new_n8911;
  assign new_n8913 = ~new_n5170 & ~new_n8912;
  assign new_n8914 = ~new_n5207 & n2184;
  assign new_n8915 = n2216 & new_n5207;
  assign new_n8916 = ~new_n8914 & ~new_n8915;
  assign new_n8917 = ~new_n5243 & ~new_n8916;
  assign new_n8918 = ~new_n5207 & n2248;
  assign new_n8919 = n2280 & new_n5207;
  assign new_n8920 = ~new_n8918 & ~new_n8919;
  assign new_n8921 = ~new_n8920 & new_n5243;
  assign new_n8922 = ~new_n8917 & ~new_n8921;
  assign new_n8923 = ~new_n8922 & new_n5170;
  assign new_n8924 = ~new_n8913 & ~new_n8923;
  assign new_n8925 = ~new_n5139 & ~new_n8924;
  assign new_n8926 = ~new_n5207 & n2312;
  assign new_n8927 = n2344 & new_n5207;
  assign new_n8928 = ~new_n8926 & ~new_n8927;
  assign new_n8929 = ~new_n5243 & ~new_n8928;
  assign new_n8930 = ~new_n5207 & n2376;
  assign new_n8931 = n2408 & new_n5207;
  assign new_n8932 = ~new_n8930 & ~new_n8931;
  assign new_n8933 = ~new_n8932 & new_n5243;
  assign new_n8934 = ~new_n8929 & ~new_n8933;
  assign new_n8935 = ~new_n5170 & ~new_n8934;
  assign new_n8936 = ~new_n5207 & n2440;
  assign new_n8937 = n2472 & new_n5207;
  assign new_n8938 = ~new_n8936 & ~new_n8937;
  assign new_n8939 = ~new_n5243 & ~new_n8938;
  assign new_n8940 = ~new_n5207 & n2504;
  assign new_n8941 = n2536 & new_n5207;
  assign new_n8942 = ~new_n8940 & ~new_n8941;
  assign new_n8943 = ~new_n8942 & new_n5243;
  assign new_n8944 = ~new_n8939 & ~new_n8943;
  assign new_n8945 = ~new_n8944 & new_n5170;
  assign new_n8946 = ~new_n8935 & ~new_n8945;
  assign new_n8947 = ~new_n8946 & new_n5139;
  assign new_n8948 = ~new_n8925 & ~new_n8947;
  assign new_n8949 = ~new_n5011 & ~new_n8948;
  assign new_n8950 = ~new_n5207 & n2568;
  assign new_n8951 = n2600 & new_n5207;
  assign new_n8952 = ~new_n8950 & ~new_n8951;
  assign new_n8953 = ~new_n5243 & ~new_n8952;
  assign new_n8954 = ~new_n5207 & n2632;
  assign new_n8955 = n2664 & new_n5207;
  assign new_n8956 = ~new_n8954 & ~new_n8955;
  assign new_n8957 = ~new_n8956 & new_n5243;
  assign new_n8958 = ~new_n8953 & ~new_n8957;
  assign new_n8959 = ~new_n5170 & ~new_n8958;
  assign new_n8960 = ~new_n5207 & n2696;
  assign new_n8961 = n2728 & new_n5207;
  assign new_n8962 = ~new_n8960 & ~new_n8961;
  assign new_n8963 = ~new_n5243 & ~new_n8962;
  assign new_n8964 = ~new_n5207 & n2760;
  assign new_n8965 = n2792 & new_n5207;
  assign new_n8966 = ~new_n8964 & ~new_n8965;
  assign new_n8967 = ~new_n8966 & new_n5243;
  assign new_n8968 = ~new_n8963 & ~new_n8967;
  assign new_n8969 = ~new_n8968 & new_n5170;
  assign new_n8970 = ~new_n8959 & ~new_n8969;
  assign new_n8971 = ~new_n5139 & ~new_n8970;
  assign new_n8972 = ~new_n5207 & n2824;
  assign new_n8973 = n2856 & new_n5207;
  assign new_n8974 = ~new_n8972 & ~new_n8973;
  assign new_n8975 = ~new_n5243 & ~new_n8974;
  assign new_n8976 = ~new_n5207 & n2888;
  assign new_n8977 = n2920 & new_n5207;
  assign new_n8978 = ~new_n8976 & ~new_n8977;
  assign new_n8979 = ~new_n8978 & new_n5243;
  assign new_n8980 = ~new_n8975 & ~new_n8979;
  assign new_n8981 = ~new_n5170 & ~new_n8980;
  assign new_n8982 = ~new_n5207 & n2952;
  assign new_n8983 = n2984 & new_n5207;
  assign new_n8984 = ~new_n8982 & ~new_n8983;
  assign new_n8985 = ~new_n5243 & ~new_n8984;
  assign new_n8986 = ~new_n5207 & n3016;
  assign new_n8987 = n3048 & new_n5207;
  assign new_n8988 = ~new_n8986 & ~new_n8987;
  assign new_n8989 = ~new_n8988 & new_n5243;
  assign new_n8990 = ~new_n8985 & ~new_n8989;
  assign new_n8991 = ~new_n8990 & new_n5170;
  assign new_n8992 = ~new_n8981 & ~new_n8991;
  assign new_n8993 = ~new_n8992 & new_n5139;
  assign new_n8994 = ~new_n8971 & ~new_n8993;
  assign new_n8995 = ~new_n8994 & new_n5011;
  assign new_n8996 = ~new_n8949 & ~new_n8995;
  assign new_n8997 = ~new_n5031 & ~new_n8996;
  assign new_n8998 = ~new_n5207 & n3080;
  assign new_n8999 = n3112 & new_n5207;
  assign new_n9000 = ~new_n8998 & ~new_n8999;
  assign new_n9001 = ~new_n5243 & ~new_n9000;
  assign new_n9002 = ~new_n5207 & n3144;
  assign new_n9003 = n3176 & new_n5207;
  assign new_n9004 = ~new_n9002 & ~new_n9003;
  assign new_n9005 = ~new_n9004 & new_n5243;
  assign new_n9006 = ~new_n9001 & ~new_n9005;
  assign new_n9007 = ~new_n5170 & ~new_n9006;
  assign new_n9008 = ~new_n5207 & n3208;
  assign new_n9009 = n3240 & new_n5207;
  assign new_n9010 = ~new_n9008 & ~new_n9009;
  assign new_n9011 = ~new_n5243 & ~new_n9010;
  assign new_n9012 = ~new_n5207 & n3272;
  assign new_n9013 = n3304 & new_n5207;
  assign new_n9014 = ~new_n9012 & ~new_n9013;
  assign new_n9015 = ~new_n9014 & new_n5243;
  assign new_n9016 = ~new_n9011 & ~new_n9015;
  assign new_n9017 = ~new_n9016 & new_n5170;
  assign new_n9018 = ~new_n9007 & ~new_n9017;
  assign new_n9019 = ~new_n5139 & ~new_n9018;
  assign new_n9020 = ~new_n5207 & n3336;
  assign new_n9021 = n3368 & new_n5207;
  assign new_n9022 = ~new_n9020 & ~new_n9021;
  assign new_n9023 = ~new_n5243 & ~new_n9022;
  assign new_n9024 = ~new_n5207 & n3400;
  assign new_n9025 = n3432 & new_n5207;
  assign new_n9026 = ~new_n9024 & ~new_n9025;
  assign new_n9027 = ~new_n9026 & new_n5243;
  assign new_n9028 = ~new_n9023 & ~new_n9027;
  assign new_n9029 = ~new_n5170 & ~new_n9028;
  assign new_n9030 = ~new_n5207 & n3464;
  assign new_n9031 = n3496 & new_n5207;
  assign new_n9032 = ~new_n9030 & ~new_n9031;
  assign new_n9033 = ~new_n5243 & ~new_n9032;
  assign new_n9034 = ~new_n5207 & n3528;
  assign new_n9035 = n3560 & new_n5207;
  assign new_n9036 = ~new_n9034 & ~new_n9035;
  assign new_n9037 = ~new_n9036 & new_n5243;
  assign new_n9038 = ~new_n9033 & ~new_n9037;
  assign new_n9039 = ~new_n9038 & new_n5170;
  assign new_n9040 = ~new_n9029 & ~new_n9039;
  assign new_n9041 = ~new_n9040 & new_n5139;
  assign new_n9042 = ~new_n9019 & ~new_n9041;
  assign new_n9043 = ~new_n5011 & ~new_n9042;
  assign new_n9044 = ~new_n5207 & n3592;
  assign new_n9045 = n3624 & new_n5207;
  assign new_n9046 = ~new_n9044 & ~new_n9045;
  assign new_n9047 = ~new_n5243 & ~new_n9046;
  assign new_n9048 = ~new_n5207 & n3656;
  assign new_n9049 = n3688 & new_n5207;
  assign new_n9050 = ~new_n9048 & ~new_n9049;
  assign new_n9051 = ~new_n9050 & new_n5243;
  assign new_n9052 = ~new_n9047 & ~new_n9051;
  assign new_n9053 = ~new_n5170 & ~new_n9052;
  assign new_n9054 = ~new_n5207 & n3720;
  assign new_n9055 = n3752 & new_n5207;
  assign new_n9056 = ~new_n9054 & ~new_n9055;
  assign new_n9057 = ~new_n5243 & ~new_n9056;
  assign new_n9058 = ~new_n5207 & n3784;
  assign new_n9059 = n3816 & new_n5207;
  assign new_n9060 = ~new_n9058 & ~new_n9059;
  assign new_n9061 = ~new_n9060 & new_n5243;
  assign new_n9062 = ~new_n9057 & ~new_n9061;
  assign new_n9063 = ~new_n9062 & new_n5170;
  assign new_n9064 = ~new_n9053 & ~new_n9063;
  assign new_n9065 = ~new_n5139 & ~new_n9064;
  assign new_n9066 = ~new_n5207 & n3848;
  assign new_n9067 = n3880 & new_n5207;
  assign new_n9068 = ~new_n9066 & ~new_n9067;
  assign new_n9069 = ~new_n5243 & ~new_n9068;
  assign new_n9070 = ~new_n5207 & n3912;
  assign new_n9071 = n3944 & new_n5207;
  assign new_n9072 = ~new_n9070 & ~new_n9071;
  assign new_n9073 = ~new_n9072 & new_n5243;
  assign new_n9074 = ~new_n9069 & ~new_n9073;
  assign new_n9075 = ~new_n5170 & ~new_n9074;
  assign new_n9076 = ~new_n5207 & n3976;
  assign new_n9077 = n4008 & new_n5207;
  assign new_n9078 = ~new_n9076 & ~new_n9077;
  assign new_n9079 = ~new_n5243 & ~new_n9078;
  assign new_n9080 = ~new_n5207 & n4040;
  assign new_n9081 = n4072 & new_n5207;
  assign new_n9082 = ~new_n9080 & ~new_n9081;
  assign new_n9083 = ~new_n9082 & new_n5243;
  assign new_n9084 = ~new_n9079 & ~new_n9083;
  assign new_n9085 = ~new_n9084 & new_n5170;
  assign new_n9086 = ~new_n9075 & ~new_n9085;
  assign new_n9087 = ~new_n9086 & new_n5139;
  assign new_n9088 = ~new_n9065 & ~new_n9087;
  assign new_n9089 = ~new_n9088 & new_n5011;
  assign new_n9090 = ~new_n9043 & ~new_n9089;
  assign new_n9091 = ~new_n9090 & new_n5031;
  assign new_n9092 = ~new_n8997 & ~new_n9091;
  assign new_n9093 = ~new_n9092 & new_n5114;
  assign new_n9094 = ~new_n5462 & ~new_n8894;
  assign new_n9095 = ~new_n9093 & ~new_n9094;
  assign new_n9096 = ~new_n5207 & n2072;
  assign new_n9097 = n2104 & new_n5207;
  assign new_n9098 = ~new_n9096 & ~new_n9097;
  assign new_n9099 = ~new_n5243 & ~new_n9098;
  assign new_n9100 = ~new_n5207 & n2136;
  assign new_n9101 = n2168 & new_n5207;
  assign new_n9102 = ~new_n9100 & ~new_n9101;
  assign new_n9103 = ~new_n9102 & new_n5243;
  assign new_n9104 = ~new_n9099 & ~new_n9103;
  assign new_n9105 = ~new_n5170 & ~new_n9104;
  assign new_n9106 = ~new_n5207 & n2200;
  assign new_n9107 = n2232 & new_n5207;
  assign new_n9108 = ~new_n9106 & ~new_n9107;
  assign new_n9109 = ~new_n5243 & ~new_n9108;
  assign new_n9110 = ~new_n5207 & n2264;
  assign new_n9111 = n2296 & new_n5207;
  assign new_n9112 = ~new_n9110 & ~new_n9111;
  assign new_n9113 = ~new_n9112 & new_n5243;
  assign new_n9114 = ~new_n9109 & ~new_n9113;
  assign new_n9115 = ~new_n9114 & new_n5170;
  assign new_n9116 = ~new_n9105 & ~new_n9115;
  assign new_n9117 = ~new_n5139 & ~new_n9116;
  assign new_n9118 = ~new_n5207 & n2328;
  assign new_n9119 = n2360 & new_n5207;
  assign new_n9120 = ~new_n9118 & ~new_n9119;
  assign new_n9121 = ~new_n5243 & ~new_n9120;
  assign new_n9122 = ~new_n5207 & n2392;
  assign new_n9123 = n2424 & new_n5207;
  assign new_n9124 = ~new_n9122 & ~new_n9123;
  assign new_n9125 = ~new_n9124 & new_n5243;
  assign new_n9126 = ~new_n9121 & ~new_n9125;
  assign new_n9127 = ~new_n5170 & ~new_n9126;
  assign new_n9128 = ~new_n5207 & n2456;
  assign new_n9129 = n2488 & new_n5207;
  assign new_n9130 = ~new_n9128 & ~new_n9129;
  assign new_n9131 = ~new_n5243 & ~new_n9130;
  assign new_n9132 = ~new_n5207 & n2520;
  assign new_n9133 = n2552 & new_n5207;
  assign new_n9134 = ~new_n9132 & ~new_n9133;
  assign new_n9135 = ~new_n9134 & new_n5243;
  assign new_n9136 = ~new_n9131 & ~new_n9135;
  assign new_n9137 = ~new_n9136 & new_n5170;
  assign new_n9138 = ~new_n9127 & ~new_n9137;
  assign new_n9139 = ~new_n9138 & new_n5139;
  assign new_n9140 = ~new_n9117 & ~new_n9139;
  assign new_n9141 = ~new_n5011 & ~new_n9140;
  assign new_n9142 = ~new_n5207 & n2584;
  assign new_n9143 = n2616 & new_n5207;
  assign new_n9144 = ~new_n9142 & ~new_n9143;
  assign new_n9145 = ~new_n5243 & ~new_n9144;
  assign new_n9146 = ~new_n5207 & n2648;
  assign new_n9147 = n2680 & new_n5207;
  assign new_n9148 = ~new_n9146 & ~new_n9147;
  assign new_n9149 = ~new_n9148 & new_n5243;
  assign new_n9150 = ~new_n9145 & ~new_n9149;
  assign new_n9151 = ~new_n5170 & ~new_n9150;
  assign new_n9152 = ~new_n5207 & n2712;
  assign new_n9153 = n2744 & new_n5207;
  assign new_n9154 = ~new_n9152 & ~new_n9153;
  assign new_n9155 = ~new_n5243 & ~new_n9154;
  assign new_n9156 = ~new_n5207 & n2776;
  assign new_n9157 = n2808 & new_n5207;
  assign new_n9158 = ~new_n9156 & ~new_n9157;
  assign new_n9159 = ~new_n9158 & new_n5243;
  assign new_n9160 = ~new_n9155 & ~new_n9159;
  assign new_n9161 = ~new_n9160 & new_n5170;
  assign new_n9162 = ~new_n9151 & ~new_n9161;
  assign new_n9163 = ~new_n5139 & ~new_n9162;
  assign new_n9164 = ~new_n5207 & n2840;
  assign new_n9165 = n2872 & new_n5207;
  assign new_n9166 = ~new_n9164 & ~new_n9165;
  assign new_n9167 = ~new_n5243 & ~new_n9166;
  assign new_n9168 = ~new_n5207 & n2904;
  assign new_n9169 = n2936 & new_n5207;
  assign new_n9170 = ~new_n9168 & ~new_n9169;
  assign new_n9171 = ~new_n9170 & new_n5243;
  assign new_n9172 = ~new_n9167 & ~new_n9171;
  assign new_n9173 = ~new_n5170 & ~new_n9172;
  assign new_n9174 = ~new_n5207 & n2968;
  assign new_n9175 = n3000 & new_n5207;
  assign new_n9176 = ~new_n9174 & ~new_n9175;
  assign new_n9177 = ~new_n5243 & ~new_n9176;
  assign new_n9178 = ~new_n5207 & n3032;
  assign new_n9179 = n3064 & new_n5207;
  assign new_n9180 = ~new_n9178 & ~new_n9179;
  assign new_n9181 = ~new_n9180 & new_n5243;
  assign new_n9182 = ~new_n9177 & ~new_n9181;
  assign new_n9183 = ~new_n9182 & new_n5170;
  assign new_n9184 = ~new_n9173 & ~new_n9183;
  assign new_n9185 = ~new_n9184 & new_n5139;
  assign new_n9186 = ~new_n9163 & ~new_n9185;
  assign new_n9187 = ~new_n9186 & new_n5011;
  assign new_n9188 = ~new_n9141 & ~new_n9187;
  assign new_n9189 = ~new_n5031 & ~new_n9188;
  assign new_n9190 = ~new_n5207 & n3096;
  assign new_n9191 = n3128 & new_n5207;
  assign new_n9192 = ~new_n9190 & ~new_n9191;
  assign new_n9193 = ~new_n5243 & ~new_n9192;
  assign new_n9194 = ~new_n5207 & n3160;
  assign new_n9195 = n3192 & new_n5207;
  assign new_n9196 = ~new_n9194 & ~new_n9195;
  assign new_n9197 = ~new_n9196 & new_n5243;
  assign new_n9198 = ~new_n9193 & ~new_n9197;
  assign new_n9199 = ~new_n5170 & ~new_n9198;
  assign new_n9200 = ~new_n5207 & n3224;
  assign new_n9201 = n3256 & new_n5207;
  assign new_n9202 = ~new_n9200 & ~new_n9201;
  assign new_n9203 = ~new_n5243 & ~new_n9202;
  assign new_n9204 = ~new_n5207 & n3288;
  assign new_n9205 = n3320 & new_n5207;
  assign new_n9206 = ~new_n9204 & ~new_n9205;
  assign new_n9207 = ~new_n9206 & new_n5243;
  assign new_n9208 = ~new_n9203 & ~new_n9207;
  assign new_n9209 = ~new_n9208 & new_n5170;
  assign new_n9210 = ~new_n9199 & ~new_n9209;
  assign new_n9211 = ~new_n5139 & ~new_n9210;
  assign new_n9212 = ~new_n5207 & n3352;
  assign new_n9213 = n3384 & new_n5207;
  assign new_n9214 = ~new_n9212 & ~new_n9213;
  assign new_n9215 = ~new_n5243 & ~new_n9214;
  assign new_n9216 = ~new_n5207 & n3416;
  assign new_n9217 = n3448 & new_n5207;
  assign new_n9218 = ~new_n9216 & ~new_n9217;
  assign new_n9219 = ~new_n9218 & new_n5243;
  assign new_n9220 = ~new_n9215 & ~new_n9219;
  assign new_n9221 = ~new_n5170 & ~new_n9220;
  assign new_n9222 = ~new_n5207 & n3480;
  assign new_n9223 = n3512 & new_n5207;
  assign new_n9224 = ~new_n9222 & ~new_n9223;
  assign new_n9225 = ~new_n5243 & ~new_n9224;
  assign new_n9226 = ~new_n5207 & n3544;
  assign new_n9227 = n3576 & new_n5207;
  assign new_n9228 = ~new_n9226 & ~new_n9227;
  assign new_n9229 = ~new_n9228 & new_n5243;
  assign new_n9230 = ~new_n9225 & ~new_n9229;
  assign new_n9231 = ~new_n9230 & new_n5170;
  assign new_n9232 = ~new_n9221 & ~new_n9231;
  assign new_n9233 = ~new_n9232 & new_n5139;
  assign new_n9234 = ~new_n9211 & ~new_n9233;
  assign new_n9235 = ~new_n5011 & ~new_n9234;
  assign new_n9236 = ~new_n5207 & n3608;
  assign new_n9237 = n3640 & new_n5207;
  assign new_n9238 = ~new_n9236 & ~new_n9237;
  assign new_n9239 = ~new_n5243 & ~new_n9238;
  assign new_n9240 = ~new_n5207 & n3672;
  assign new_n9241 = n3704 & new_n5207;
  assign new_n9242 = ~new_n9240 & ~new_n9241;
  assign new_n9243 = ~new_n9242 & new_n5243;
  assign new_n9244 = ~new_n9239 & ~new_n9243;
  assign new_n9245 = ~new_n5170 & ~new_n9244;
  assign new_n9246 = ~new_n5207 & n3736;
  assign new_n9247 = n3768 & new_n5207;
  assign new_n9248 = ~new_n9246 & ~new_n9247;
  assign new_n9249 = ~new_n5243 & ~new_n9248;
  assign new_n9250 = ~new_n5207 & n3800;
  assign new_n9251 = n3832 & new_n5207;
  assign new_n9252 = ~new_n9250 & ~new_n9251;
  assign new_n9253 = ~new_n9252 & new_n5243;
  assign new_n9254 = ~new_n9249 & ~new_n9253;
  assign new_n9255 = ~new_n9254 & new_n5170;
  assign new_n9256 = ~new_n9245 & ~new_n9255;
  assign new_n9257 = ~new_n5139 & ~new_n9256;
  assign new_n9258 = ~new_n5207 & n3864;
  assign new_n9259 = n3896 & new_n5207;
  assign new_n9260 = ~new_n9258 & ~new_n9259;
  assign new_n9261 = ~new_n5243 & ~new_n9260;
  assign new_n9262 = ~new_n5207 & n3928;
  assign new_n9263 = n3960 & new_n5207;
  assign new_n9264 = ~new_n9262 & ~new_n9263;
  assign new_n9265 = ~new_n9264 & new_n5243;
  assign new_n9266 = ~new_n9261 & ~new_n9265;
  assign new_n9267 = ~new_n5170 & ~new_n9266;
  assign new_n9268 = ~new_n5207 & n3992;
  assign new_n9269 = n4024 & new_n5207;
  assign new_n9270 = ~new_n9268 & ~new_n9269;
  assign new_n9271 = ~new_n5243 & ~new_n9270;
  assign new_n9272 = ~new_n5207 & n4056;
  assign new_n9273 = n4088 & new_n5207;
  assign new_n9274 = ~new_n9272 & ~new_n9273;
  assign new_n9275 = ~new_n9274 & new_n5243;
  assign new_n9276 = ~new_n9271 & ~new_n9275;
  assign new_n9277 = ~new_n9276 & new_n5170;
  assign new_n9278 = ~new_n9267 & ~new_n9277;
  assign new_n9279 = ~new_n9278 & new_n5139;
  assign new_n9280 = ~new_n9257 & ~new_n9279;
  assign new_n9281 = ~new_n9280 & new_n5011;
  assign new_n9282 = ~new_n9235 & ~new_n9281;
  assign new_n9283 = ~new_n9282 & new_n5031;
  assign new_n9284 = ~new_n9189 & ~new_n9283;
  assign new_n9285 = ~new_n5115 & ~new_n9284;
  assign new_n9286 = ~new_n5116 & ~new_n8704;
  assign new_n9287 = ~new_n9285 & ~new_n9286;
  assign new_n9288 = new_n9095 & new_n9287;
  assign new_n9289 = new_n8900 ^ new_n8899;
  assign new_n9290 = ~new_n9288 & ~new_n9289;
  assign new_n9291 = ~new_n8903 & ~new_n9290;
  assign new_n9292 = ~new_n4113 & new_n4270;
  assign new_n9293 = ~new_n4107 & ~new_n9292;
  assign new_n9294 = new_n8421 ^ new_n4106;
  assign new_n9295 = ~new_n9293 & ~new_n9294;
  assign new_n9296 = new_n9295 ^ new_n4260;
  assign new_n9297 = ~new_n9296 & new_n4118;
  assign new_n9298 = new_n4117 ^ n2019;
  assign new_n9299 = ~new_n9297 & ~new_n9298;
  assign new_n9300 = ~new_n4129 & ~new_n4137;
  assign new_n9301 = new_n9299 & new_n9300;
  assign new_n9302 = new_n9301 ^ new_n4138;
  assign new_n9303 = ~new_n5113 & ~new_n9302;
  assign new_n9304 = ~new_n9303 & new_n9291;
  assign new_n9305 = ~new_n8896 & new_n8901;
  assign new_n9306 = ~new_n8704 & new_n4150;
  assign new_n9307 = ~new_n9305 & ~new_n9306;
  assign new_n9308 = ~new_n9288 & new_n8900;
  assign new_n9309 = ~new_n9308 & new_n9307;
  assign new_n9310 = new_n9304 & new_n9309;
  assign new_n9311 = ~new_n9310 & new_n8515;
  assign new_n9312 = ~new_n5207 & n2063;
  assign new_n9313 = n2095 & new_n5207;
  assign new_n9314 = ~new_n9312 & ~new_n9313;
  assign new_n9315 = ~new_n5243 & ~new_n9314;
  assign new_n9316 = ~new_n5207 & n2127;
  assign new_n9317 = n2159 & new_n5207;
  assign new_n9318 = ~new_n9316 & ~new_n9317;
  assign new_n9319 = ~new_n9318 & new_n5243;
  assign new_n9320 = ~new_n9315 & ~new_n9319;
  assign new_n9321 = ~new_n5170 & ~new_n9320;
  assign new_n9322 = ~new_n5207 & n2191;
  assign new_n9323 = n2223 & new_n5207;
  assign new_n9324 = ~new_n9322 & ~new_n9323;
  assign new_n9325 = ~new_n5243 & ~new_n9324;
  assign new_n9326 = ~new_n5207 & n2255;
  assign new_n9327 = n2287 & new_n5207;
  assign new_n9328 = ~new_n9326 & ~new_n9327;
  assign new_n9329 = ~new_n9328 & new_n5243;
  assign new_n9330 = ~new_n9325 & ~new_n9329;
  assign new_n9331 = ~new_n9330 & new_n5170;
  assign new_n9332 = ~new_n9321 & ~new_n9331;
  assign new_n9333 = ~new_n5139 & ~new_n9332;
  assign new_n9334 = ~new_n5207 & n2319;
  assign new_n9335 = n2351 & new_n5207;
  assign new_n9336 = ~new_n9334 & ~new_n9335;
  assign new_n9337 = ~new_n5243 & ~new_n9336;
  assign new_n9338 = ~new_n5207 & n2383;
  assign new_n9339 = n2415 & new_n5207;
  assign new_n9340 = ~new_n9338 & ~new_n9339;
  assign new_n9341 = ~new_n9340 & new_n5243;
  assign new_n9342 = ~new_n9337 & ~new_n9341;
  assign new_n9343 = ~new_n5170 & ~new_n9342;
  assign new_n9344 = ~new_n5207 & n2447;
  assign new_n9345 = n2479 & new_n5207;
  assign new_n9346 = ~new_n9344 & ~new_n9345;
  assign new_n9347 = ~new_n5243 & ~new_n9346;
  assign new_n9348 = ~new_n5207 & n2511;
  assign new_n9349 = n2543 & new_n5207;
  assign new_n9350 = ~new_n9348 & ~new_n9349;
  assign new_n9351 = ~new_n9350 & new_n5243;
  assign new_n9352 = ~new_n9347 & ~new_n9351;
  assign new_n9353 = ~new_n9352 & new_n5170;
  assign new_n9354 = ~new_n9343 & ~new_n9353;
  assign new_n9355 = ~new_n9354 & new_n5139;
  assign new_n9356 = ~new_n9333 & ~new_n9355;
  assign new_n9357 = ~new_n5011 & ~new_n9356;
  assign new_n9358 = ~new_n5207 & n2575;
  assign new_n9359 = n2607 & new_n5207;
  assign new_n9360 = ~new_n9358 & ~new_n9359;
  assign new_n9361 = ~new_n5243 & ~new_n9360;
  assign new_n9362 = ~new_n5207 & n2639;
  assign new_n9363 = n2671 & new_n5207;
  assign new_n9364 = ~new_n9362 & ~new_n9363;
  assign new_n9365 = ~new_n9364 & new_n5243;
  assign new_n9366 = ~new_n9361 & ~new_n9365;
  assign new_n9367 = ~new_n5170 & ~new_n9366;
  assign new_n9368 = ~new_n5207 & n2703;
  assign new_n9369 = n2735 & new_n5207;
  assign new_n9370 = ~new_n9368 & ~new_n9369;
  assign new_n9371 = ~new_n5243 & ~new_n9370;
  assign new_n9372 = ~new_n5207 & n2767;
  assign new_n9373 = n2799 & new_n5207;
  assign new_n9374 = ~new_n9372 & ~new_n9373;
  assign new_n9375 = ~new_n9374 & new_n5243;
  assign new_n9376 = ~new_n9371 & ~new_n9375;
  assign new_n9377 = ~new_n9376 & new_n5170;
  assign new_n9378 = ~new_n9367 & ~new_n9377;
  assign new_n9379 = ~new_n5139 & ~new_n9378;
  assign new_n9380 = ~new_n5207 & n2831;
  assign new_n9381 = n2863 & new_n5207;
  assign new_n9382 = ~new_n9380 & ~new_n9381;
  assign new_n9383 = ~new_n5243 & ~new_n9382;
  assign new_n9384 = ~new_n5207 & n2895;
  assign new_n9385 = n2927 & new_n5207;
  assign new_n9386 = ~new_n9384 & ~new_n9385;
  assign new_n9387 = ~new_n9386 & new_n5243;
  assign new_n9388 = ~new_n9383 & ~new_n9387;
  assign new_n9389 = ~new_n5170 & ~new_n9388;
  assign new_n9390 = ~new_n5207 & n2959;
  assign new_n9391 = n2991 & new_n5207;
  assign new_n9392 = ~new_n9390 & ~new_n9391;
  assign new_n9393 = ~new_n5243 & ~new_n9392;
  assign new_n9394 = ~new_n5207 & n3023;
  assign new_n9395 = n3055 & new_n5207;
  assign new_n9396 = ~new_n9394 & ~new_n9395;
  assign new_n9397 = ~new_n9396 & new_n5243;
  assign new_n9398 = ~new_n9393 & ~new_n9397;
  assign new_n9399 = ~new_n9398 & new_n5170;
  assign new_n9400 = ~new_n9389 & ~new_n9399;
  assign new_n9401 = ~new_n9400 & new_n5139;
  assign new_n9402 = ~new_n9379 & ~new_n9401;
  assign new_n9403 = ~new_n9402 & new_n5011;
  assign new_n9404 = ~new_n9357 & ~new_n9403;
  assign new_n9405 = ~new_n5031 & ~new_n9404;
  assign new_n9406 = ~new_n5207 & n3087;
  assign new_n9407 = n3119 & new_n5207;
  assign new_n9408 = ~new_n9406 & ~new_n9407;
  assign new_n9409 = ~new_n5243 & ~new_n9408;
  assign new_n9410 = ~new_n5207 & n3151;
  assign new_n9411 = n3183 & new_n5207;
  assign new_n9412 = ~new_n9410 & ~new_n9411;
  assign new_n9413 = ~new_n9412 & new_n5243;
  assign new_n9414 = ~new_n9409 & ~new_n9413;
  assign new_n9415 = ~new_n5170 & ~new_n9414;
  assign new_n9416 = ~new_n5207 & n3215;
  assign new_n9417 = n3247 & new_n5207;
  assign new_n9418 = ~new_n9416 & ~new_n9417;
  assign new_n9419 = ~new_n5243 & ~new_n9418;
  assign new_n9420 = ~new_n5207 & n3279;
  assign new_n9421 = n3311 & new_n5207;
  assign new_n9422 = ~new_n9420 & ~new_n9421;
  assign new_n9423 = ~new_n9422 & new_n5243;
  assign new_n9424 = ~new_n9419 & ~new_n9423;
  assign new_n9425 = ~new_n9424 & new_n5170;
  assign new_n9426 = ~new_n9415 & ~new_n9425;
  assign new_n9427 = ~new_n5139 & ~new_n9426;
  assign new_n9428 = ~new_n5207 & n3343;
  assign new_n9429 = n3375 & new_n5207;
  assign new_n9430 = ~new_n9428 & ~new_n9429;
  assign new_n9431 = ~new_n5243 & ~new_n9430;
  assign new_n9432 = ~new_n5207 & n3407;
  assign new_n9433 = n3439 & new_n5207;
  assign new_n9434 = ~new_n9432 & ~new_n9433;
  assign new_n9435 = ~new_n9434 & new_n5243;
  assign new_n9436 = ~new_n9431 & ~new_n9435;
  assign new_n9437 = ~new_n5170 & ~new_n9436;
  assign new_n9438 = ~new_n5207 & n3471;
  assign new_n9439 = n3503 & new_n5207;
  assign new_n9440 = ~new_n9438 & ~new_n9439;
  assign new_n9441 = ~new_n5243 & ~new_n9440;
  assign new_n9442 = ~new_n5207 & n3535;
  assign new_n9443 = n3567 & new_n5207;
  assign new_n9444 = ~new_n9442 & ~new_n9443;
  assign new_n9445 = ~new_n9444 & new_n5243;
  assign new_n9446 = ~new_n9441 & ~new_n9445;
  assign new_n9447 = ~new_n9446 & new_n5170;
  assign new_n9448 = ~new_n9437 & ~new_n9447;
  assign new_n9449 = ~new_n9448 & new_n5139;
  assign new_n9450 = ~new_n9427 & ~new_n9449;
  assign new_n9451 = ~new_n5011 & ~new_n9450;
  assign new_n9452 = ~new_n5207 & n3599;
  assign new_n9453 = n3631 & new_n5207;
  assign new_n9454 = ~new_n9452 & ~new_n9453;
  assign new_n9455 = ~new_n5243 & ~new_n9454;
  assign new_n9456 = ~new_n5207 & n3663;
  assign new_n9457 = n3695 & new_n5207;
  assign new_n9458 = ~new_n9456 & ~new_n9457;
  assign new_n9459 = ~new_n9458 & new_n5243;
  assign new_n9460 = ~new_n9455 & ~new_n9459;
  assign new_n9461 = ~new_n5170 & ~new_n9460;
  assign new_n9462 = ~new_n5207 & n3727;
  assign new_n9463 = n3759 & new_n5207;
  assign new_n9464 = ~new_n9462 & ~new_n9463;
  assign new_n9465 = ~new_n5243 & ~new_n9464;
  assign new_n9466 = ~new_n5207 & n3791;
  assign new_n9467 = n3823 & new_n5207;
  assign new_n9468 = ~new_n9466 & ~new_n9467;
  assign new_n9469 = ~new_n9468 & new_n5243;
  assign new_n9470 = ~new_n9465 & ~new_n9469;
  assign new_n9471 = ~new_n9470 & new_n5170;
  assign new_n9472 = ~new_n9461 & ~new_n9471;
  assign new_n9473 = ~new_n5139 & ~new_n9472;
  assign new_n9474 = ~new_n5207 & n3855;
  assign new_n9475 = n3887 & new_n5207;
  assign new_n9476 = ~new_n9474 & ~new_n9475;
  assign new_n9477 = ~new_n5243 & ~new_n9476;
  assign new_n9478 = ~new_n5207 & n3919;
  assign new_n9479 = n3951 & new_n5207;
  assign new_n9480 = ~new_n9478 & ~new_n9479;
  assign new_n9481 = ~new_n9480 & new_n5243;
  assign new_n9482 = ~new_n9477 & ~new_n9481;
  assign new_n9483 = ~new_n5170 & ~new_n9482;
  assign new_n9484 = ~new_n5207 & n3983;
  assign new_n9485 = n4015 & new_n5207;
  assign new_n9486 = ~new_n9484 & ~new_n9485;
  assign new_n9487 = ~new_n5243 & ~new_n9486;
  assign new_n9488 = ~new_n5207 & n4047;
  assign new_n9489 = n4079 & new_n5207;
  assign new_n9490 = ~new_n9488 & ~new_n9489;
  assign new_n9491 = ~new_n9490 & new_n5243;
  assign new_n9492 = ~new_n9487 & ~new_n9491;
  assign new_n9493 = ~new_n9492 & new_n5170;
  assign new_n9494 = ~new_n9483 & ~new_n9493;
  assign new_n9495 = ~new_n9494 & new_n5139;
  assign new_n9496 = ~new_n9473 & ~new_n9495;
  assign new_n9497 = ~new_n9496 & new_n5011;
  assign new_n9498 = ~new_n9451 & ~new_n9497;
  assign new_n9499 = ~new_n9498 & new_n5031;
  assign new_n9500 = ~new_n9405 & ~new_n9499;
  assign new_n9501 = ~new_n5077 & ~new_n9500;
  assign new_n9502 = ~new_n5207 & n2079;
  assign new_n9503 = n2111 & new_n5207;
  assign new_n9504 = ~new_n9502 & ~new_n9503;
  assign new_n9505 = ~new_n5243 & ~new_n9504;
  assign new_n9506 = ~new_n5207 & n2143;
  assign new_n9507 = n2175 & new_n5207;
  assign new_n9508 = ~new_n9506 & ~new_n9507;
  assign new_n9509 = ~new_n9508 & new_n5243;
  assign new_n9510 = ~new_n9505 & ~new_n9509;
  assign new_n9511 = ~new_n5170 & ~new_n9510;
  assign new_n9512 = ~new_n5207 & n2207;
  assign new_n9513 = n2239 & new_n5207;
  assign new_n9514 = ~new_n9512 & ~new_n9513;
  assign new_n9515 = ~new_n5243 & ~new_n9514;
  assign new_n9516 = ~new_n5207 & n2271;
  assign new_n9517 = n2303 & new_n5207;
  assign new_n9518 = ~new_n9516 & ~new_n9517;
  assign new_n9519 = ~new_n9518 & new_n5243;
  assign new_n9520 = ~new_n9515 & ~new_n9519;
  assign new_n9521 = ~new_n9520 & new_n5170;
  assign new_n9522 = ~new_n9511 & ~new_n9521;
  assign new_n9523 = ~new_n5139 & ~new_n9522;
  assign new_n9524 = ~new_n5207 & n2335;
  assign new_n9525 = n2367 & new_n5207;
  assign new_n9526 = ~new_n9524 & ~new_n9525;
  assign new_n9527 = ~new_n5243 & ~new_n9526;
  assign new_n9528 = ~new_n5207 & n2399;
  assign new_n9529 = n2431 & new_n5207;
  assign new_n9530 = ~new_n9528 & ~new_n9529;
  assign new_n9531 = ~new_n9530 & new_n5243;
  assign new_n9532 = ~new_n9527 & ~new_n9531;
  assign new_n9533 = ~new_n5170 & ~new_n9532;
  assign new_n9534 = ~new_n5207 & n2463;
  assign new_n9535 = n2495 & new_n5207;
  assign new_n9536 = ~new_n9534 & ~new_n9535;
  assign new_n9537 = ~new_n5243 & ~new_n9536;
  assign new_n9538 = ~new_n5207 & n2527;
  assign new_n9539 = n2559 & new_n5207;
  assign new_n9540 = ~new_n9538 & ~new_n9539;
  assign new_n9541 = ~new_n9540 & new_n5243;
  assign new_n9542 = ~new_n9537 & ~new_n9541;
  assign new_n9543 = ~new_n9542 & new_n5170;
  assign new_n9544 = ~new_n9533 & ~new_n9543;
  assign new_n9545 = ~new_n9544 & new_n5139;
  assign new_n9546 = ~new_n9523 & ~new_n9545;
  assign new_n9547 = ~new_n5011 & ~new_n9546;
  assign new_n9548 = ~new_n5207 & n2591;
  assign new_n9549 = n2623 & new_n5207;
  assign new_n9550 = ~new_n9548 & ~new_n9549;
  assign new_n9551 = ~new_n5243 & ~new_n9550;
  assign new_n9552 = ~new_n5207 & n2655;
  assign new_n9553 = n2687 & new_n5207;
  assign new_n9554 = ~new_n9552 & ~new_n9553;
  assign new_n9555 = ~new_n9554 & new_n5243;
  assign new_n9556 = ~new_n9551 & ~new_n9555;
  assign new_n9557 = ~new_n5170 & ~new_n9556;
  assign new_n9558 = ~new_n5207 & n2719;
  assign new_n9559 = n2751 & new_n5207;
  assign new_n9560 = ~new_n9558 & ~new_n9559;
  assign new_n9561 = ~new_n5243 & ~new_n9560;
  assign new_n9562 = ~new_n5207 & n2783;
  assign new_n9563 = n2815 & new_n5207;
  assign new_n9564 = ~new_n9562 & ~new_n9563;
  assign new_n9565 = ~new_n9564 & new_n5243;
  assign new_n9566 = ~new_n9561 & ~new_n9565;
  assign new_n9567 = ~new_n9566 & new_n5170;
  assign new_n9568 = ~new_n9557 & ~new_n9567;
  assign new_n9569 = ~new_n5139 & ~new_n9568;
  assign new_n9570 = ~new_n5207 & n2847;
  assign new_n9571 = n2879 & new_n5207;
  assign new_n9572 = ~new_n9570 & ~new_n9571;
  assign new_n9573 = ~new_n5243 & ~new_n9572;
  assign new_n9574 = ~new_n5207 & n2911;
  assign new_n9575 = n2943 & new_n5207;
  assign new_n9576 = ~new_n9574 & ~new_n9575;
  assign new_n9577 = ~new_n9576 & new_n5243;
  assign new_n9578 = ~new_n9573 & ~new_n9577;
  assign new_n9579 = ~new_n5170 & ~new_n9578;
  assign new_n9580 = ~new_n5207 & n2975;
  assign new_n9581 = n3007 & new_n5207;
  assign new_n9582 = ~new_n9580 & ~new_n9581;
  assign new_n9583 = ~new_n5243 & ~new_n9582;
  assign new_n9584 = ~new_n5207 & n3039;
  assign new_n9585 = n3071 & new_n5207;
  assign new_n9586 = ~new_n9584 & ~new_n9585;
  assign new_n9587 = ~new_n9586 & new_n5243;
  assign new_n9588 = ~new_n9583 & ~new_n9587;
  assign new_n9589 = ~new_n9588 & new_n5170;
  assign new_n9590 = ~new_n9579 & ~new_n9589;
  assign new_n9591 = ~new_n9590 & new_n5139;
  assign new_n9592 = ~new_n9569 & ~new_n9591;
  assign new_n9593 = ~new_n9592 & new_n5011;
  assign new_n9594 = ~new_n9547 & ~new_n9593;
  assign new_n9595 = ~new_n5031 & ~new_n9594;
  assign new_n9596 = ~new_n5207 & n3103;
  assign new_n9597 = n3135 & new_n5207;
  assign new_n9598 = ~new_n9596 & ~new_n9597;
  assign new_n9599 = ~new_n5243 & ~new_n9598;
  assign new_n9600 = ~new_n5207 & n3167;
  assign new_n9601 = n3199 & new_n5207;
  assign new_n9602 = ~new_n9600 & ~new_n9601;
  assign new_n9603 = ~new_n9602 & new_n5243;
  assign new_n9604 = ~new_n9599 & ~new_n9603;
  assign new_n9605 = ~new_n5170 & ~new_n9604;
  assign new_n9606 = ~new_n5207 & n3231;
  assign new_n9607 = n3263 & new_n5207;
  assign new_n9608 = ~new_n9606 & ~new_n9607;
  assign new_n9609 = ~new_n5243 & ~new_n9608;
  assign new_n9610 = ~new_n5207 & n3295;
  assign new_n9611 = n3327 & new_n5207;
  assign new_n9612 = ~new_n9610 & ~new_n9611;
  assign new_n9613 = ~new_n9612 & new_n5243;
  assign new_n9614 = ~new_n9609 & ~new_n9613;
  assign new_n9615 = ~new_n9614 & new_n5170;
  assign new_n9616 = ~new_n9605 & ~new_n9615;
  assign new_n9617 = ~new_n5139 & ~new_n9616;
  assign new_n9618 = ~new_n5207 & n3359;
  assign new_n9619 = n3391 & new_n5207;
  assign new_n9620 = ~new_n9618 & ~new_n9619;
  assign new_n9621 = ~new_n5243 & ~new_n9620;
  assign new_n9622 = ~new_n5207 & n3423;
  assign new_n9623 = n3455 & new_n5207;
  assign new_n9624 = ~new_n9622 & ~new_n9623;
  assign new_n9625 = ~new_n9624 & new_n5243;
  assign new_n9626 = ~new_n9621 & ~new_n9625;
  assign new_n9627 = ~new_n5170 & ~new_n9626;
  assign new_n9628 = ~new_n5207 & n3487;
  assign new_n9629 = n3519 & new_n5207;
  assign new_n9630 = ~new_n9628 & ~new_n9629;
  assign new_n9631 = ~new_n5243 & ~new_n9630;
  assign new_n9632 = ~new_n5207 & n3551;
  assign new_n9633 = n3583 & new_n5207;
  assign new_n9634 = ~new_n9632 & ~new_n9633;
  assign new_n9635 = ~new_n9634 & new_n5243;
  assign new_n9636 = ~new_n9631 & ~new_n9635;
  assign new_n9637 = ~new_n9636 & new_n5170;
  assign new_n9638 = ~new_n9627 & ~new_n9637;
  assign new_n9639 = ~new_n9638 & new_n5139;
  assign new_n9640 = ~new_n9617 & ~new_n9639;
  assign new_n9641 = ~new_n5011 & ~new_n9640;
  assign new_n9642 = ~new_n5207 & n3615;
  assign new_n9643 = n3647 & new_n5207;
  assign new_n9644 = ~new_n9642 & ~new_n9643;
  assign new_n9645 = ~new_n5243 & ~new_n9644;
  assign new_n9646 = ~new_n5207 & n3679;
  assign new_n9647 = n3711 & new_n5207;
  assign new_n9648 = ~new_n9646 & ~new_n9647;
  assign new_n9649 = ~new_n9648 & new_n5243;
  assign new_n9650 = ~new_n9645 & ~new_n9649;
  assign new_n9651 = ~new_n5170 & ~new_n9650;
  assign new_n9652 = ~new_n5207 & n3743;
  assign new_n9653 = n3775 & new_n5207;
  assign new_n9654 = ~new_n9652 & ~new_n9653;
  assign new_n9655 = ~new_n5243 & ~new_n9654;
  assign new_n9656 = ~new_n5207 & n3807;
  assign new_n9657 = n3839 & new_n5207;
  assign new_n9658 = ~new_n9656 & ~new_n9657;
  assign new_n9659 = ~new_n9658 & new_n5243;
  assign new_n9660 = ~new_n9655 & ~new_n9659;
  assign new_n9661 = ~new_n9660 & new_n5170;
  assign new_n9662 = ~new_n9651 & ~new_n9661;
  assign new_n9663 = ~new_n5139 & ~new_n9662;
  assign new_n9664 = ~new_n5207 & n3871;
  assign new_n9665 = n3903 & new_n5207;
  assign new_n9666 = ~new_n9664 & ~new_n9665;
  assign new_n9667 = ~new_n5243 & ~new_n9666;
  assign new_n9668 = ~new_n5207 & n3935;
  assign new_n9669 = n3967 & new_n5207;
  assign new_n9670 = ~new_n9668 & ~new_n9669;
  assign new_n9671 = ~new_n9670 & new_n5243;
  assign new_n9672 = ~new_n9667 & ~new_n9671;
  assign new_n9673 = ~new_n5170 & ~new_n9672;
  assign new_n9674 = ~new_n5207 & n3999;
  assign new_n9675 = n4031 & new_n5207;
  assign new_n9676 = ~new_n9674 & ~new_n9675;
  assign new_n9677 = ~new_n5243 & ~new_n9676;
  assign new_n9678 = ~new_n5207 & n4063;
  assign new_n9679 = n4095 & new_n5207;
  assign new_n9680 = ~new_n9678 & ~new_n9679;
  assign new_n9681 = ~new_n9680 & new_n5243;
  assign new_n9682 = ~new_n9677 & ~new_n9681;
  assign new_n9683 = ~new_n9682 & new_n5170;
  assign new_n9684 = ~new_n9673 & ~new_n9683;
  assign new_n9685 = ~new_n9684 & new_n5139;
  assign new_n9686 = ~new_n9663 & ~new_n9685;
  assign new_n9687 = ~new_n9686 & new_n5011;
  assign new_n9688 = ~new_n9641 & ~new_n9687;
  assign new_n9689 = ~new_n9688 & new_n5031;
  assign new_n9690 = ~new_n9595 & ~new_n9689;
  assign new_n9691 = ~new_n9690 & new_n5077;
  assign new_n9692 = ~new_n9501 & ~new_n9691;
  assign new_n9693 = ~new_n9692 & new_n8902;
  assign new_n9694 = ~new_n5207 & n2055;
  assign new_n9695 = n2087 & new_n5207;
  assign new_n9696 = ~new_n9694 & ~new_n9695;
  assign new_n9697 = ~new_n5243 & ~new_n9696;
  assign new_n9698 = ~new_n5207 & n2119;
  assign new_n9699 = n2151 & new_n5207;
  assign new_n9700 = ~new_n9698 & ~new_n9699;
  assign new_n9701 = ~new_n9700 & new_n5243;
  assign new_n9702 = ~new_n9697 & ~new_n9701;
  assign new_n9703 = ~new_n5170 & ~new_n9702;
  assign new_n9704 = ~new_n5207 & n2183;
  assign new_n9705 = n2215 & new_n5207;
  assign new_n9706 = ~new_n9704 & ~new_n9705;
  assign new_n9707 = ~new_n5243 & ~new_n9706;
  assign new_n9708 = ~new_n5207 & n2247;
  assign new_n9709 = n2279 & new_n5207;
  assign new_n9710 = ~new_n9708 & ~new_n9709;
  assign new_n9711 = ~new_n9710 & new_n5243;
  assign new_n9712 = ~new_n9707 & ~new_n9711;
  assign new_n9713 = ~new_n9712 & new_n5170;
  assign new_n9714 = ~new_n9703 & ~new_n9713;
  assign new_n9715 = ~new_n5139 & ~new_n9714;
  assign new_n9716 = ~new_n5207 & n2311;
  assign new_n9717 = n2343 & new_n5207;
  assign new_n9718 = ~new_n9716 & ~new_n9717;
  assign new_n9719 = ~new_n5243 & ~new_n9718;
  assign new_n9720 = ~new_n5207 & n2375;
  assign new_n9721 = n2407 & new_n5207;
  assign new_n9722 = ~new_n9720 & ~new_n9721;
  assign new_n9723 = ~new_n9722 & new_n5243;
  assign new_n9724 = ~new_n9719 & ~new_n9723;
  assign new_n9725 = ~new_n5170 & ~new_n9724;
  assign new_n9726 = ~new_n5207 & n2439;
  assign new_n9727 = n2471 & new_n5207;
  assign new_n9728 = ~new_n9726 & ~new_n9727;
  assign new_n9729 = ~new_n5243 & ~new_n9728;
  assign new_n9730 = ~new_n5207 & n2503;
  assign new_n9731 = n2535 & new_n5207;
  assign new_n9732 = ~new_n9730 & ~new_n9731;
  assign new_n9733 = ~new_n9732 & new_n5243;
  assign new_n9734 = ~new_n9729 & ~new_n9733;
  assign new_n9735 = ~new_n9734 & new_n5170;
  assign new_n9736 = ~new_n9725 & ~new_n9735;
  assign new_n9737 = ~new_n9736 & new_n5139;
  assign new_n9738 = ~new_n9715 & ~new_n9737;
  assign new_n9739 = ~new_n5011 & ~new_n9738;
  assign new_n9740 = ~new_n5207 & n2567;
  assign new_n9741 = n2599 & new_n5207;
  assign new_n9742 = ~new_n9740 & ~new_n9741;
  assign new_n9743 = ~new_n5243 & ~new_n9742;
  assign new_n9744 = ~new_n5207 & n2631;
  assign new_n9745 = n2663 & new_n5207;
  assign new_n9746 = ~new_n9744 & ~new_n9745;
  assign new_n9747 = ~new_n9746 & new_n5243;
  assign new_n9748 = ~new_n9743 & ~new_n9747;
  assign new_n9749 = ~new_n5170 & ~new_n9748;
  assign new_n9750 = ~new_n5207 & n2695;
  assign new_n9751 = n2727 & new_n5207;
  assign new_n9752 = ~new_n9750 & ~new_n9751;
  assign new_n9753 = ~new_n5243 & ~new_n9752;
  assign new_n9754 = ~new_n5207 & n2759;
  assign new_n9755 = n2791 & new_n5207;
  assign new_n9756 = ~new_n9754 & ~new_n9755;
  assign new_n9757 = ~new_n9756 & new_n5243;
  assign new_n9758 = ~new_n9753 & ~new_n9757;
  assign new_n9759 = ~new_n9758 & new_n5170;
  assign new_n9760 = ~new_n9749 & ~new_n9759;
  assign new_n9761 = ~new_n5139 & ~new_n9760;
  assign new_n9762 = ~new_n5207 & n2823;
  assign new_n9763 = n2855 & new_n5207;
  assign new_n9764 = ~new_n9762 & ~new_n9763;
  assign new_n9765 = ~new_n5243 & ~new_n9764;
  assign new_n9766 = ~new_n5207 & n2887;
  assign new_n9767 = n2919 & new_n5207;
  assign new_n9768 = ~new_n9766 & ~new_n9767;
  assign new_n9769 = ~new_n9768 & new_n5243;
  assign new_n9770 = ~new_n9765 & ~new_n9769;
  assign new_n9771 = ~new_n5170 & ~new_n9770;
  assign new_n9772 = ~new_n5207 & n2951;
  assign new_n9773 = n2983 & new_n5207;
  assign new_n9774 = ~new_n9772 & ~new_n9773;
  assign new_n9775 = ~new_n5243 & ~new_n9774;
  assign new_n9776 = ~new_n5207 & n3015;
  assign new_n9777 = n3047 & new_n5207;
  assign new_n9778 = ~new_n9776 & ~new_n9777;
  assign new_n9779 = ~new_n9778 & new_n5243;
  assign new_n9780 = ~new_n9775 & ~new_n9779;
  assign new_n9781 = ~new_n9780 & new_n5170;
  assign new_n9782 = ~new_n9771 & ~new_n9781;
  assign new_n9783 = ~new_n9782 & new_n5139;
  assign new_n9784 = ~new_n9761 & ~new_n9783;
  assign new_n9785 = ~new_n9784 & new_n5011;
  assign new_n9786 = ~new_n9739 & ~new_n9785;
  assign new_n9787 = ~new_n5031 & ~new_n9786;
  assign new_n9788 = ~new_n5207 & n3079;
  assign new_n9789 = n3111 & new_n5207;
  assign new_n9790 = ~new_n9788 & ~new_n9789;
  assign new_n9791 = ~new_n5243 & ~new_n9790;
  assign new_n9792 = ~new_n5207 & n3143;
  assign new_n9793 = n3175 & new_n5207;
  assign new_n9794 = ~new_n9792 & ~new_n9793;
  assign new_n9795 = ~new_n9794 & new_n5243;
  assign new_n9796 = ~new_n9791 & ~new_n9795;
  assign new_n9797 = ~new_n5170 & ~new_n9796;
  assign new_n9798 = ~new_n5207 & n3207;
  assign new_n9799 = n3239 & new_n5207;
  assign new_n9800 = ~new_n9798 & ~new_n9799;
  assign new_n9801 = ~new_n5243 & ~new_n9800;
  assign new_n9802 = ~new_n5207 & n3271;
  assign new_n9803 = n3303 & new_n5207;
  assign new_n9804 = ~new_n9802 & ~new_n9803;
  assign new_n9805 = ~new_n9804 & new_n5243;
  assign new_n9806 = ~new_n9801 & ~new_n9805;
  assign new_n9807 = ~new_n9806 & new_n5170;
  assign new_n9808 = ~new_n9797 & ~new_n9807;
  assign new_n9809 = ~new_n5139 & ~new_n9808;
  assign new_n9810 = ~new_n5207 & n3335;
  assign new_n9811 = n3367 & new_n5207;
  assign new_n9812 = ~new_n9810 & ~new_n9811;
  assign new_n9813 = ~new_n5243 & ~new_n9812;
  assign new_n9814 = ~new_n5207 & n3399;
  assign new_n9815 = n3431 & new_n5207;
  assign new_n9816 = ~new_n9814 & ~new_n9815;
  assign new_n9817 = ~new_n9816 & new_n5243;
  assign new_n9818 = ~new_n9813 & ~new_n9817;
  assign new_n9819 = ~new_n5170 & ~new_n9818;
  assign new_n9820 = ~new_n5207 & n3463;
  assign new_n9821 = n3495 & new_n5207;
  assign new_n9822 = ~new_n9820 & ~new_n9821;
  assign new_n9823 = ~new_n5243 & ~new_n9822;
  assign new_n9824 = ~new_n5207 & n3527;
  assign new_n9825 = n3559 & new_n5207;
  assign new_n9826 = ~new_n9824 & ~new_n9825;
  assign new_n9827 = ~new_n9826 & new_n5243;
  assign new_n9828 = ~new_n9823 & ~new_n9827;
  assign new_n9829 = ~new_n9828 & new_n5170;
  assign new_n9830 = ~new_n9819 & ~new_n9829;
  assign new_n9831 = ~new_n9830 & new_n5139;
  assign new_n9832 = ~new_n9809 & ~new_n9831;
  assign new_n9833 = ~new_n5011 & ~new_n9832;
  assign new_n9834 = ~new_n5207 & n3591;
  assign new_n9835 = n3623 & new_n5207;
  assign new_n9836 = ~new_n9834 & ~new_n9835;
  assign new_n9837 = ~new_n5243 & ~new_n9836;
  assign new_n9838 = ~new_n5207 & n3655;
  assign new_n9839 = n3687 & new_n5207;
  assign new_n9840 = ~new_n9838 & ~new_n9839;
  assign new_n9841 = ~new_n9840 & new_n5243;
  assign new_n9842 = ~new_n9837 & ~new_n9841;
  assign new_n9843 = ~new_n5170 & ~new_n9842;
  assign new_n9844 = ~new_n5207 & n3719;
  assign new_n9845 = n3751 & new_n5207;
  assign new_n9846 = ~new_n9844 & ~new_n9845;
  assign new_n9847 = ~new_n5243 & ~new_n9846;
  assign new_n9848 = ~new_n5207 & n3783;
  assign new_n9849 = n3815 & new_n5207;
  assign new_n9850 = ~new_n9848 & ~new_n9849;
  assign new_n9851 = ~new_n9850 & new_n5243;
  assign new_n9852 = ~new_n9847 & ~new_n9851;
  assign new_n9853 = ~new_n9852 & new_n5170;
  assign new_n9854 = ~new_n9843 & ~new_n9853;
  assign new_n9855 = ~new_n5139 & ~new_n9854;
  assign new_n9856 = ~new_n5207 & n3847;
  assign new_n9857 = n3879 & new_n5207;
  assign new_n9858 = ~new_n9856 & ~new_n9857;
  assign new_n9859 = ~new_n5243 & ~new_n9858;
  assign new_n9860 = ~new_n5207 & n3911;
  assign new_n9861 = n3943 & new_n5207;
  assign new_n9862 = ~new_n9860 & ~new_n9861;
  assign new_n9863 = ~new_n9862 & new_n5243;
  assign new_n9864 = ~new_n9859 & ~new_n9863;
  assign new_n9865 = ~new_n5170 & ~new_n9864;
  assign new_n9866 = ~new_n5207 & n3975;
  assign new_n9867 = n4007 & new_n5207;
  assign new_n9868 = ~new_n9866 & ~new_n9867;
  assign new_n9869 = ~new_n5243 & ~new_n9868;
  assign new_n9870 = ~new_n5207 & n4039;
  assign new_n9871 = n4071 & new_n5207;
  assign new_n9872 = ~new_n9870 & ~new_n9871;
  assign new_n9873 = ~new_n9872 & new_n5243;
  assign new_n9874 = ~new_n9869 & ~new_n9873;
  assign new_n9875 = ~new_n9874 & new_n5170;
  assign new_n9876 = ~new_n9865 & ~new_n9875;
  assign new_n9877 = ~new_n9876 & new_n5139;
  assign new_n9878 = ~new_n9855 & ~new_n9877;
  assign new_n9879 = ~new_n9878 & new_n5011;
  assign new_n9880 = ~new_n9833 & ~new_n9879;
  assign new_n9881 = ~new_n9880 & new_n5031;
  assign new_n9882 = ~new_n9787 & ~new_n9881;
  assign new_n9883 = ~new_n9882 & new_n5114;
  assign new_n9884 = ~new_n5462 & ~new_n9500;
  assign new_n9885 = ~new_n9883 & ~new_n9884;
  assign new_n9886 = ~new_n5207 & n2071;
  assign new_n9887 = n2103 & new_n5207;
  assign new_n9888 = ~new_n9886 & ~new_n9887;
  assign new_n9889 = ~new_n5243 & ~new_n9888;
  assign new_n9890 = ~new_n5207 & n2135;
  assign new_n9891 = n2167 & new_n5207;
  assign new_n9892 = ~new_n9890 & ~new_n9891;
  assign new_n9893 = ~new_n9892 & new_n5243;
  assign new_n9894 = ~new_n9889 & ~new_n9893;
  assign new_n9895 = ~new_n5170 & ~new_n9894;
  assign new_n9896 = ~new_n5207 & n2199;
  assign new_n9897 = n2231 & new_n5207;
  assign new_n9898 = ~new_n9896 & ~new_n9897;
  assign new_n9899 = ~new_n5243 & ~new_n9898;
  assign new_n9900 = ~new_n5207 & n2263;
  assign new_n9901 = n2295 & new_n5207;
  assign new_n9902 = ~new_n9900 & ~new_n9901;
  assign new_n9903 = ~new_n9902 & new_n5243;
  assign new_n9904 = ~new_n9899 & ~new_n9903;
  assign new_n9905 = ~new_n9904 & new_n5170;
  assign new_n9906 = ~new_n9895 & ~new_n9905;
  assign new_n9907 = ~new_n5139 & ~new_n9906;
  assign new_n9908 = ~new_n5207 & n2327;
  assign new_n9909 = n2359 & new_n5207;
  assign new_n9910 = ~new_n9908 & ~new_n9909;
  assign new_n9911 = ~new_n5243 & ~new_n9910;
  assign new_n9912 = ~new_n5207 & n2391;
  assign new_n9913 = n2423 & new_n5207;
  assign new_n9914 = ~new_n9912 & ~new_n9913;
  assign new_n9915 = ~new_n9914 & new_n5243;
  assign new_n9916 = ~new_n9911 & ~new_n9915;
  assign new_n9917 = ~new_n5170 & ~new_n9916;
  assign new_n9918 = ~new_n5207 & n2455;
  assign new_n9919 = n2487 & new_n5207;
  assign new_n9920 = ~new_n9918 & ~new_n9919;
  assign new_n9921 = ~new_n5243 & ~new_n9920;
  assign new_n9922 = ~new_n5207 & n2519;
  assign new_n9923 = n2551 & new_n5207;
  assign new_n9924 = ~new_n9922 & ~new_n9923;
  assign new_n9925 = ~new_n9924 & new_n5243;
  assign new_n9926 = ~new_n9921 & ~new_n9925;
  assign new_n9927 = ~new_n9926 & new_n5170;
  assign new_n9928 = ~new_n9917 & ~new_n9927;
  assign new_n9929 = ~new_n9928 & new_n5139;
  assign new_n9930 = ~new_n9907 & ~new_n9929;
  assign new_n9931 = ~new_n5011 & ~new_n9930;
  assign new_n9932 = ~new_n5207 & n2583;
  assign new_n9933 = n2615 & new_n5207;
  assign new_n9934 = ~new_n9932 & ~new_n9933;
  assign new_n9935 = ~new_n5243 & ~new_n9934;
  assign new_n9936 = ~new_n5207 & n2647;
  assign new_n9937 = n2679 & new_n5207;
  assign new_n9938 = ~new_n9936 & ~new_n9937;
  assign new_n9939 = ~new_n9938 & new_n5243;
  assign new_n9940 = ~new_n9935 & ~new_n9939;
  assign new_n9941 = ~new_n5170 & ~new_n9940;
  assign new_n9942 = ~new_n5207 & n2711;
  assign new_n9943 = n2743 & new_n5207;
  assign new_n9944 = ~new_n9942 & ~new_n9943;
  assign new_n9945 = ~new_n5243 & ~new_n9944;
  assign new_n9946 = ~new_n5207 & n2775;
  assign new_n9947 = n2807 & new_n5207;
  assign new_n9948 = ~new_n9946 & ~new_n9947;
  assign new_n9949 = ~new_n9948 & new_n5243;
  assign new_n9950 = ~new_n9945 & ~new_n9949;
  assign new_n9951 = ~new_n9950 & new_n5170;
  assign new_n9952 = ~new_n9941 & ~new_n9951;
  assign new_n9953 = ~new_n5139 & ~new_n9952;
  assign new_n9954 = ~new_n5207 & n2839;
  assign new_n9955 = n2871 & new_n5207;
  assign new_n9956 = ~new_n9954 & ~new_n9955;
  assign new_n9957 = ~new_n5243 & ~new_n9956;
  assign new_n9958 = ~new_n5207 & n2903;
  assign new_n9959 = n2935 & new_n5207;
  assign new_n9960 = ~new_n9958 & ~new_n9959;
  assign new_n9961 = ~new_n9960 & new_n5243;
  assign new_n9962 = ~new_n9957 & ~new_n9961;
  assign new_n9963 = ~new_n5170 & ~new_n9962;
  assign new_n9964 = ~new_n5207 & n2967;
  assign new_n9965 = n2999 & new_n5207;
  assign new_n9966 = ~new_n9964 & ~new_n9965;
  assign new_n9967 = ~new_n5243 & ~new_n9966;
  assign new_n9968 = ~new_n5207 & n3031;
  assign new_n9969 = n3063 & new_n5207;
  assign new_n9970 = ~new_n9968 & ~new_n9969;
  assign new_n9971 = ~new_n9970 & new_n5243;
  assign new_n9972 = ~new_n9967 & ~new_n9971;
  assign new_n9973 = ~new_n9972 & new_n5170;
  assign new_n9974 = ~new_n9963 & ~new_n9973;
  assign new_n9975 = ~new_n9974 & new_n5139;
  assign new_n9976 = ~new_n9953 & ~new_n9975;
  assign new_n9977 = ~new_n9976 & new_n5011;
  assign new_n9978 = ~new_n9931 & ~new_n9977;
  assign new_n9979 = ~new_n5031 & ~new_n9978;
  assign new_n9980 = ~new_n5207 & n3095;
  assign new_n9981 = n3127 & new_n5207;
  assign new_n9982 = ~new_n9980 & ~new_n9981;
  assign new_n9983 = ~new_n5243 & ~new_n9982;
  assign new_n9984 = ~new_n5207 & n3159;
  assign new_n9985 = n3191 & new_n5207;
  assign new_n9986 = ~new_n9984 & ~new_n9985;
  assign new_n9987 = ~new_n9986 & new_n5243;
  assign new_n9988 = ~new_n9983 & ~new_n9987;
  assign new_n9989 = ~new_n5170 & ~new_n9988;
  assign new_n9990 = ~new_n5207 & n3223;
  assign new_n9991 = n3255 & new_n5207;
  assign new_n9992 = ~new_n9990 & ~new_n9991;
  assign new_n9993 = ~new_n5243 & ~new_n9992;
  assign new_n9994 = ~new_n5207 & n3287;
  assign new_n9995 = n3319 & new_n5207;
  assign new_n9996 = ~new_n9994 & ~new_n9995;
  assign new_n9997 = ~new_n9996 & new_n5243;
  assign new_n9998 = ~new_n9993 & ~new_n9997;
  assign new_n9999 = ~new_n9998 & new_n5170;
  assign new_n10000 = ~new_n9989 & ~new_n9999;
  assign new_n10001 = ~new_n5139 & ~new_n10000;
  assign new_n10002 = ~new_n5207 & n3351;
  assign new_n10003 = n3383 & new_n5207;
  assign new_n10004 = ~new_n10002 & ~new_n10003;
  assign new_n10005 = ~new_n5243 & ~new_n10004;
  assign new_n10006 = ~new_n5207 & n3415;
  assign new_n10007 = n3447 & new_n5207;
  assign new_n10008 = ~new_n10006 & ~new_n10007;
  assign new_n10009 = ~new_n10008 & new_n5243;
  assign new_n10010 = ~new_n10005 & ~new_n10009;
  assign new_n10011 = ~new_n5170 & ~new_n10010;
  assign new_n10012 = ~new_n5207 & n3479;
  assign new_n10013 = n3511 & new_n5207;
  assign new_n10014 = ~new_n10012 & ~new_n10013;
  assign new_n10015 = ~new_n5243 & ~new_n10014;
  assign new_n10016 = ~new_n5207 & n3543;
  assign new_n10017 = n3575 & new_n5207;
  assign new_n10018 = ~new_n10016 & ~new_n10017;
  assign new_n10019 = ~new_n10018 & new_n5243;
  assign new_n10020 = ~new_n10015 & ~new_n10019;
  assign new_n10021 = ~new_n10020 & new_n5170;
  assign new_n10022 = ~new_n10011 & ~new_n10021;
  assign new_n10023 = ~new_n10022 & new_n5139;
  assign new_n10024 = ~new_n10001 & ~new_n10023;
  assign new_n10025 = ~new_n5011 & ~new_n10024;
  assign new_n10026 = ~new_n5207 & n3607;
  assign new_n10027 = n3639 & new_n5207;
  assign new_n10028 = ~new_n10026 & ~new_n10027;
  assign new_n10029 = ~new_n5243 & ~new_n10028;
  assign new_n10030 = ~new_n5207 & n3671;
  assign new_n10031 = n3703 & new_n5207;
  assign new_n10032 = ~new_n10030 & ~new_n10031;
  assign new_n10033 = ~new_n10032 & new_n5243;
  assign new_n10034 = ~new_n10029 & ~new_n10033;
  assign new_n10035 = ~new_n5170 & ~new_n10034;
  assign new_n10036 = ~new_n5207 & n3735;
  assign new_n10037 = n3767 & new_n5207;
  assign new_n10038 = ~new_n10036 & ~new_n10037;
  assign new_n10039 = ~new_n5243 & ~new_n10038;
  assign new_n10040 = ~new_n5207 & n3799;
  assign new_n10041 = n3831 & new_n5207;
  assign new_n10042 = ~new_n10040 & ~new_n10041;
  assign new_n10043 = ~new_n10042 & new_n5243;
  assign new_n10044 = ~new_n10039 & ~new_n10043;
  assign new_n10045 = ~new_n10044 & new_n5170;
  assign new_n10046 = ~new_n10035 & ~new_n10045;
  assign new_n10047 = ~new_n5139 & ~new_n10046;
  assign new_n10048 = ~new_n5207 & n3863;
  assign new_n10049 = n3895 & new_n5207;
  assign new_n10050 = ~new_n10048 & ~new_n10049;
  assign new_n10051 = ~new_n5243 & ~new_n10050;
  assign new_n10052 = ~new_n5207 & n3927;
  assign new_n10053 = n3959 & new_n5207;
  assign new_n10054 = ~new_n10052 & ~new_n10053;
  assign new_n10055 = ~new_n10054 & new_n5243;
  assign new_n10056 = ~new_n10051 & ~new_n10055;
  assign new_n10057 = ~new_n5170 & ~new_n10056;
  assign new_n10058 = ~new_n5207 & n3991;
  assign new_n10059 = n4023 & new_n5207;
  assign new_n10060 = ~new_n10058 & ~new_n10059;
  assign new_n10061 = ~new_n5243 & ~new_n10060;
  assign new_n10062 = ~new_n5207 & n4055;
  assign new_n10063 = n4087 & new_n5207;
  assign new_n10064 = ~new_n10062 & ~new_n10063;
  assign new_n10065 = ~new_n10064 & new_n5243;
  assign new_n10066 = ~new_n10061 & ~new_n10065;
  assign new_n10067 = ~new_n10066 & new_n5170;
  assign new_n10068 = ~new_n10057 & ~new_n10067;
  assign new_n10069 = ~new_n10068 & new_n5139;
  assign new_n10070 = ~new_n10047 & ~new_n10069;
  assign new_n10071 = ~new_n10070 & new_n5011;
  assign new_n10072 = ~new_n10025 & ~new_n10071;
  assign new_n10073 = ~new_n10072 & new_n5031;
  assign new_n10074 = ~new_n9979 & ~new_n10073;
  assign new_n10075 = ~new_n5115 & ~new_n10074;
  assign new_n10076 = ~new_n5116 & ~new_n9690;
  assign new_n10077 = ~new_n10075 & ~new_n10076;
  assign new_n10078 = new_n9885 & new_n10077;
  assign new_n10079 = ~new_n9289 & ~new_n10078;
  assign new_n10080 = ~new_n9693 & ~new_n10079;
  assign new_n10081 = ~new_n5077 & ~new_n9302;
  assign new_n10082 = ~new_n10081 & new_n10080;
  assign new_n10083 = ~new_n9692 & new_n8901;
  assign new_n10084 = ~new_n9690 & new_n4150;
  assign new_n10085 = ~new_n10083 & ~new_n10084;
  assign new_n10086 = ~new_n10078 & new_n8900;
  assign new_n10087 = ~new_n10086 & new_n10085;
  assign new_n10088 = new_n10082 & new_n10087;
  assign new_n10089 = ~new_n10088 & new_n8515;
  assign new_n10090 = new_n4135 ^ n2020;
  assign new_n10091 = new_n10090 ^ new_n9295;
  assign new_n10092 = new_n4118 & new_n10091;
  assign new_n10093 = ~new_n5207 & n2062;
  assign new_n10094 = n2094 & new_n5207;
  assign new_n10095 = ~new_n10093 & ~new_n10094;
  assign new_n10096 = ~new_n5243 & ~new_n10095;
  assign new_n10097 = ~new_n5207 & n2126;
  assign new_n10098 = n2158 & new_n5207;
  assign new_n10099 = ~new_n10097 & ~new_n10098;
  assign new_n10100 = ~new_n10099 & new_n5243;
  assign new_n10101 = ~new_n10096 & ~new_n10100;
  assign new_n10102 = ~new_n5170 & ~new_n10101;
  assign new_n10103 = ~new_n5207 & n2190;
  assign new_n10104 = n2222 & new_n5207;
  assign new_n10105 = ~new_n10103 & ~new_n10104;
  assign new_n10106 = ~new_n5243 & ~new_n10105;
  assign new_n10107 = ~new_n5207 & n2254;
  assign new_n10108 = n2286 & new_n5207;
  assign new_n10109 = ~new_n10107 & ~new_n10108;
  assign new_n10110 = ~new_n10109 & new_n5243;
  assign new_n10111 = ~new_n10106 & ~new_n10110;
  assign new_n10112 = ~new_n10111 & new_n5170;
  assign new_n10113 = ~new_n10102 & ~new_n10112;
  assign new_n10114 = ~new_n5139 & ~new_n10113;
  assign new_n10115 = ~new_n5207 & n2318;
  assign new_n10116 = n2350 & new_n5207;
  assign new_n10117 = ~new_n10115 & ~new_n10116;
  assign new_n10118 = ~new_n5243 & ~new_n10117;
  assign new_n10119 = ~new_n5207 & n2382;
  assign new_n10120 = n2414 & new_n5207;
  assign new_n10121 = ~new_n10119 & ~new_n10120;
  assign new_n10122 = ~new_n10121 & new_n5243;
  assign new_n10123 = ~new_n10118 & ~new_n10122;
  assign new_n10124 = ~new_n5170 & ~new_n10123;
  assign new_n10125 = ~new_n5207 & n2446;
  assign new_n10126 = n2478 & new_n5207;
  assign new_n10127 = ~new_n10125 & ~new_n10126;
  assign new_n10128 = ~new_n5243 & ~new_n10127;
  assign new_n10129 = ~new_n5207 & n2510;
  assign new_n10130 = n2542 & new_n5207;
  assign new_n10131 = ~new_n10129 & ~new_n10130;
  assign new_n10132 = ~new_n10131 & new_n5243;
  assign new_n10133 = ~new_n10128 & ~new_n10132;
  assign new_n10134 = ~new_n10133 & new_n5170;
  assign new_n10135 = ~new_n10124 & ~new_n10134;
  assign new_n10136 = ~new_n10135 & new_n5139;
  assign new_n10137 = ~new_n10114 & ~new_n10136;
  assign new_n10138 = ~new_n5011 & ~new_n10137;
  assign new_n10139 = ~new_n5207 & n2574;
  assign new_n10140 = n2606 & new_n5207;
  assign new_n10141 = ~new_n10139 & ~new_n10140;
  assign new_n10142 = ~new_n5243 & ~new_n10141;
  assign new_n10143 = ~new_n5207 & n2638;
  assign new_n10144 = n2670 & new_n5207;
  assign new_n10145 = ~new_n10143 & ~new_n10144;
  assign new_n10146 = ~new_n10145 & new_n5243;
  assign new_n10147 = ~new_n10142 & ~new_n10146;
  assign new_n10148 = ~new_n5170 & ~new_n10147;
  assign new_n10149 = ~new_n5207 & n2702;
  assign new_n10150 = n2734 & new_n5207;
  assign new_n10151 = ~new_n10149 & ~new_n10150;
  assign new_n10152 = ~new_n5243 & ~new_n10151;
  assign new_n10153 = ~new_n5207 & n2766;
  assign new_n10154 = n2798 & new_n5207;
  assign new_n10155 = ~new_n10153 & ~new_n10154;
  assign new_n10156 = ~new_n10155 & new_n5243;
  assign new_n10157 = ~new_n10152 & ~new_n10156;
  assign new_n10158 = ~new_n10157 & new_n5170;
  assign new_n10159 = ~new_n10148 & ~new_n10158;
  assign new_n10160 = ~new_n5139 & ~new_n10159;
  assign new_n10161 = ~new_n5207 & n2830;
  assign new_n10162 = n2862 & new_n5207;
  assign new_n10163 = ~new_n10161 & ~new_n10162;
  assign new_n10164 = ~new_n5243 & ~new_n10163;
  assign new_n10165 = ~new_n5207 & n2894;
  assign new_n10166 = n2926 & new_n5207;
  assign new_n10167 = ~new_n10165 & ~new_n10166;
  assign new_n10168 = ~new_n10167 & new_n5243;
  assign new_n10169 = ~new_n10164 & ~new_n10168;
  assign new_n10170 = ~new_n5170 & ~new_n10169;
  assign new_n10171 = ~new_n5207 & n2958;
  assign new_n10172 = n2990 & new_n5207;
  assign new_n10173 = ~new_n10171 & ~new_n10172;
  assign new_n10174 = ~new_n5243 & ~new_n10173;
  assign new_n10175 = ~new_n5207 & n3022;
  assign new_n10176 = n3054 & new_n5207;
  assign new_n10177 = ~new_n10175 & ~new_n10176;
  assign new_n10178 = ~new_n10177 & new_n5243;
  assign new_n10179 = ~new_n10174 & ~new_n10178;
  assign new_n10180 = ~new_n10179 & new_n5170;
  assign new_n10181 = ~new_n10170 & ~new_n10180;
  assign new_n10182 = ~new_n10181 & new_n5139;
  assign new_n10183 = ~new_n10160 & ~new_n10182;
  assign new_n10184 = ~new_n10183 & new_n5011;
  assign new_n10185 = ~new_n10138 & ~new_n10184;
  assign new_n10186 = ~new_n5031 & ~new_n10185;
  assign new_n10187 = ~new_n5207 & n3086;
  assign new_n10188 = n3118 & new_n5207;
  assign new_n10189 = ~new_n10187 & ~new_n10188;
  assign new_n10190 = ~new_n5243 & ~new_n10189;
  assign new_n10191 = ~new_n5207 & n3150;
  assign new_n10192 = n3182 & new_n5207;
  assign new_n10193 = ~new_n10191 & ~new_n10192;
  assign new_n10194 = ~new_n10193 & new_n5243;
  assign new_n10195 = ~new_n10190 & ~new_n10194;
  assign new_n10196 = ~new_n5170 & ~new_n10195;
  assign new_n10197 = ~new_n5207 & n3214;
  assign new_n10198 = n3246 & new_n5207;
  assign new_n10199 = ~new_n10197 & ~new_n10198;
  assign new_n10200 = ~new_n5243 & ~new_n10199;
  assign new_n10201 = ~new_n5207 & n3278;
  assign new_n10202 = n3310 & new_n5207;
  assign new_n10203 = ~new_n10201 & ~new_n10202;
  assign new_n10204 = ~new_n10203 & new_n5243;
  assign new_n10205 = ~new_n10200 & ~new_n10204;
  assign new_n10206 = ~new_n10205 & new_n5170;
  assign new_n10207 = ~new_n10196 & ~new_n10206;
  assign new_n10208 = ~new_n5139 & ~new_n10207;
  assign new_n10209 = ~new_n5207 & n3342;
  assign new_n10210 = n3374 & new_n5207;
  assign new_n10211 = ~new_n10209 & ~new_n10210;
  assign new_n10212 = ~new_n5243 & ~new_n10211;
  assign new_n10213 = ~new_n5207 & n3406;
  assign new_n10214 = n3438 & new_n5207;
  assign new_n10215 = ~new_n10213 & ~new_n10214;
  assign new_n10216 = ~new_n10215 & new_n5243;
  assign new_n10217 = ~new_n10212 & ~new_n10216;
  assign new_n10218 = ~new_n5170 & ~new_n10217;
  assign new_n10219 = ~new_n5207 & n3470;
  assign new_n10220 = n3502 & new_n5207;
  assign new_n10221 = ~new_n10219 & ~new_n10220;
  assign new_n10222 = ~new_n5243 & ~new_n10221;
  assign new_n10223 = ~new_n5207 & n3534;
  assign new_n10224 = n3566 & new_n5207;
  assign new_n10225 = ~new_n10223 & ~new_n10224;
  assign new_n10226 = ~new_n10225 & new_n5243;
  assign new_n10227 = ~new_n10222 & ~new_n10226;
  assign new_n10228 = ~new_n10227 & new_n5170;
  assign new_n10229 = ~new_n10218 & ~new_n10228;
  assign new_n10230 = ~new_n10229 & new_n5139;
  assign new_n10231 = ~new_n10208 & ~new_n10230;
  assign new_n10232 = ~new_n5011 & ~new_n10231;
  assign new_n10233 = ~new_n5207 & n3598;
  assign new_n10234 = n3630 & new_n5207;
  assign new_n10235 = ~new_n10233 & ~new_n10234;
  assign new_n10236 = ~new_n5243 & ~new_n10235;
  assign new_n10237 = ~new_n5207 & n3662;
  assign new_n10238 = n3694 & new_n5207;
  assign new_n10239 = ~new_n10237 & ~new_n10238;
  assign new_n10240 = ~new_n10239 & new_n5243;
  assign new_n10241 = ~new_n10236 & ~new_n10240;
  assign new_n10242 = ~new_n5170 & ~new_n10241;
  assign new_n10243 = ~new_n5207 & n3726;
  assign new_n10244 = n3758 & new_n5207;
  assign new_n10245 = ~new_n10243 & ~new_n10244;
  assign new_n10246 = ~new_n5243 & ~new_n10245;
  assign new_n10247 = ~new_n5207 & n3790;
  assign new_n10248 = n3822 & new_n5207;
  assign new_n10249 = ~new_n10247 & ~new_n10248;
  assign new_n10250 = ~new_n10249 & new_n5243;
  assign new_n10251 = ~new_n10246 & ~new_n10250;
  assign new_n10252 = ~new_n10251 & new_n5170;
  assign new_n10253 = ~new_n10242 & ~new_n10252;
  assign new_n10254 = ~new_n5139 & ~new_n10253;
  assign new_n10255 = ~new_n5207 & n3854;
  assign new_n10256 = n3886 & new_n5207;
  assign new_n10257 = ~new_n10255 & ~new_n10256;
  assign new_n10258 = ~new_n5243 & ~new_n10257;
  assign new_n10259 = ~new_n5207 & n3918;
  assign new_n10260 = n3950 & new_n5207;
  assign new_n10261 = ~new_n10259 & ~new_n10260;
  assign new_n10262 = ~new_n10261 & new_n5243;
  assign new_n10263 = ~new_n10258 & ~new_n10262;
  assign new_n10264 = ~new_n5170 & ~new_n10263;
  assign new_n10265 = ~new_n5207 & n3982;
  assign new_n10266 = n4014 & new_n5207;
  assign new_n10267 = ~new_n10265 & ~new_n10266;
  assign new_n10268 = ~new_n5243 & ~new_n10267;
  assign new_n10269 = ~new_n5207 & n4046;
  assign new_n10270 = n4078 & new_n5207;
  assign new_n10271 = ~new_n10269 & ~new_n10270;
  assign new_n10272 = ~new_n10271 & new_n5243;
  assign new_n10273 = ~new_n10268 & ~new_n10272;
  assign new_n10274 = ~new_n10273 & new_n5170;
  assign new_n10275 = ~new_n10264 & ~new_n10274;
  assign new_n10276 = ~new_n10275 & new_n5139;
  assign new_n10277 = ~new_n10254 & ~new_n10276;
  assign new_n10278 = ~new_n10277 & new_n5011;
  assign new_n10279 = ~new_n10232 & ~new_n10278;
  assign new_n10280 = ~new_n10279 & new_n5031;
  assign new_n10281 = ~new_n10186 & ~new_n10280;
  assign new_n10282 = ~new_n5077 & ~new_n10281;
  assign new_n10283 = ~new_n5207 & n2078;
  assign new_n10284 = n2110 & new_n5207;
  assign new_n10285 = ~new_n10283 & ~new_n10284;
  assign new_n10286 = ~new_n5243 & ~new_n10285;
  assign new_n10287 = ~new_n5207 & n2142;
  assign new_n10288 = n2174 & new_n5207;
  assign new_n10289 = ~new_n10287 & ~new_n10288;
  assign new_n10290 = ~new_n10289 & new_n5243;
  assign new_n10291 = ~new_n10286 & ~new_n10290;
  assign new_n10292 = ~new_n5170 & ~new_n10291;
  assign new_n10293 = ~new_n5207 & n2206;
  assign new_n10294 = n2238 & new_n5207;
  assign new_n10295 = ~new_n10293 & ~new_n10294;
  assign new_n10296 = ~new_n5243 & ~new_n10295;
  assign new_n10297 = ~new_n5207 & n2270;
  assign new_n10298 = n2302 & new_n5207;
  assign new_n10299 = ~new_n10297 & ~new_n10298;
  assign new_n10300 = ~new_n10299 & new_n5243;
  assign new_n10301 = ~new_n10296 & ~new_n10300;
  assign new_n10302 = ~new_n10301 & new_n5170;
  assign new_n10303 = ~new_n10292 & ~new_n10302;
  assign new_n10304 = ~new_n5139 & ~new_n10303;
  assign new_n10305 = ~new_n5207 & n2334;
  assign new_n10306 = n2366 & new_n5207;
  assign new_n10307 = ~new_n10305 & ~new_n10306;
  assign new_n10308 = ~new_n5243 & ~new_n10307;
  assign new_n10309 = ~new_n5207 & n2398;
  assign new_n10310 = n2430 & new_n5207;
  assign new_n10311 = ~new_n10309 & ~new_n10310;
  assign new_n10312 = ~new_n10311 & new_n5243;
  assign new_n10313 = ~new_n10308 & ~new_n10312;
  assign new_n10314 = ~new_n5170 & ~new_n10313;
  assign new_n10315 = ~new_n5207 & n2462;
  assign new_n10316 = n2494 & new_n5207;
  assign new_n10317 = ~new_n10315 & ~new_n10316;
  assign new_n10318 = ~new_n5243 & ~new_n10317;
  assign new_n10319 = ~new_n5207 & n2526;
  assign new_n10320 = n2558 & new_n5207;
  assign new_n10321 = ~new_n10319 & ~new_n10320;
  assign new_n10322 = ~new_n10321 & new_n5243;
  assign new_n10323 = ~new_n10318 & ~new_n10322;
  assign new_n10324 = ~new_n10323 & new_n5170;
  assign new_n10325 = ~new_n10314 & ~new_n10324;
  assign new_n10326 = ~new_n10325 & new_n5139;
  assign new_n10327 = ~new_n10304 & ~new_n10326;
  assign new_n10328 = ~new_n5011 & ~new_n10327;
  assign new_n10329 = ~new_n5207 & n2590;
  assign new_n10330 = n2622 & new_n5207;
  assign new_n10331 = ~new_n10329 & ~new_n10330;
  assign new_n10332 = ~new_n5243 & ~new_n10331;
  assign new_n10333 = ~new_n5207 & n2654;
  assign new_n10334 = n2686 & new_n5207;
  assign new_n10335 = ~new_n10333 & ~new_n10334;
  assign new_n10336 = ~new_n10335 & new_n5243;
  assign new_n10337 = ~new_n10332 & ~new_n10336;
  assign new_n10338 = ~new_n5170 & ~new_n10337;
  assign new_n10339 = ~new_n5207 & n2718;
  assign new_n10340 = n2750 & new_n5207;
  assign new_n10341 = ~new_n10339 & ~new_n10340;
  assign new_n10342 = ~new_n5243 & ~new_n10341;
  assign new_n10343 = ~new_n5207 & n2782;
  assign new_n10344 = n2814 & new_n5207;
  assign new_n10345 = ~new_n10343 & ~new_n10344;
  assign new_n10346 = ~new_n10345 & new_n5243;
  assign new_n10347 = ~new_n10342 & ~new_n10346;
  assign new_n10348 = ~new_n10347 & new_n5170;
  assign new_n10349 = ~new_n10338 & ~new_n10348;
  assign new_n10350 = ~new_n5139 & ~new_n10349;
  assign new_n10351 = ~new_n5207 & n2846;
  assign new_n10352 = n2878 & new_n5207;
  assign new_n10353 = ~new_n10351 & ~new_n10352;
  assign new_n10354 = ~new_n5243 & ~new_n10353;
  assign new_n10355 = ~new_n5207 & n2910;
  assign new_n10356 = n2942 & new_n5207;
  assign new_n10357 = ~new_n10355 & ~new_n10356;
  assign new_n10358 = ~new_n10357 & new_n5243;
  assign new_n10359 = ~new_n10354 & ~new_n10358;
  assign new_n10360 = ~new_n5170 & ~new_n10359;
  assign new_n10361 = ~new_n5207 & n2974;
  assign new_n10362 = n3006 & new_n5207;
  assign new_n10363 = ~new_n10361 & ~new_n10362;
  assign new_n10364 = ~new_n5243 & ~new_n10363;
  assign new_n10365 = ~new_n5207 & n3038;
  assign new_n10366 = n3070 & new_n5207;
  assign new_n10367 = ~new_n10365 & ~new_n10366;
  assign new_n10368 = ~new_n10367 & new_n5243;
  assign new_n10369 = ~new_n10364 & ~new_n10368;
  assign new_n10370 = ~new_n10369 & new_n5170;
  assign new_n10371 = ~new_n10360 & ~new_n10370;
  assign new_n10372 = ~new_n10371 & new_n5139;
  assign new_n10373 = ~new_n10350 & ~new_n10372;
  assign new_n10374 = ~new_n10373 & new_n5011;
  assign new_n10375 = ~new_n10328 & ~new_n10374;
  assign new_n10376 = ~new_n5031 & ~new_n10375;
  assign new_n10377 = ~new_n5207 & n3102;
  assign new_n10378 = n3134 & new_n5207;
  assign new_n10379 = ~new_n10377 & ~new_n10378;
  assign new_n10380 = ~new_n5243 & ~new_n10379;
  assign new_n10381 = ~new_n5207 & n3166;
  assign new_n10382 = n3198 & new_n5207;
  assign new_n10383 = ~new_n10381 & ~new_n10382;
  assign new_n10384 = ~new_n10383 & new_n5243;
  assign new_n10385 = ~new_n10380 & ~new_n10384;
  assign new_n10386 = ~new_n5170 & ~new_n10385;
  assign new_n10387 = ~new_n5207 & n3230;
  assign new_n10388 = n3262 & new_n5207;
  assign new_n10389 = ~new_n10387 & ~new_n10388;
  assign new_n10390 = ~new_n5243 & ~new_n10389;
  assign new_n10391 = ~new_n5207 & n3294;
  assign new_n10392 = n3326 & new_n5207;
  assign new_n10393 = ~new_n10391 & ~new_n10392;
  assign new_n10394 = ~new_n10393 & new_n5243;
  assign new_n10395 = ~new_n10390 & ~new_n10394;
  assign new_n10396 = ~new_n10395 & new_n5170;
  assign new_n10397 = ~new_n10386 & ~new_n10396;
  assign new_n10398 = ~new_n5139 & ~new_n10397;
  assign new_n10399 = ~new_n5207 & n3358;
  assign new_n10400 = n3390 & new_n5207;
  assign new_n10401 = ~new_n10399 & ~new_n10400;
  assign new_n10402 = ~new_n5243 & ~new_n10401;
  assign new_n10403 = ~new_n5207 & n3422;
  assign new_n10404 = n3454 & new_n5207;
  assign new_n10405 = ~new_n10403 & ~new_n10404;
  assign new_n10406 = ~new_n10405 & new_n5243;
  assign new_n10407 = ~new_n10402 & ~new_n10406;
  assign new_n10408 = ~new_n5170 & ~new_n10407;
  assign new_n10409 = ~new_n5207 & n3486;
  assign new_n10410 = n3518 & new_n5207;
  assign new_n10411 = ~new_n10409 & ~new_n10410;
  assign new_n10412 = ~new_n5243 & ~new_n10411;
  assign new_n10413 = ~new_n5207 & n3550;
  assign new_n10414 = n3582 & new_n5207;
  assign new_n10415 = ~new_n10413 & ~new_n10414;
  assign new_n10416 = ~new_n10415 & new_n5243;
  assign new_n10417 = ~new_n10412 & ~new_n10416;
  assign new_n10418 = ~new_n10417 & new_n5170;
  assign new_n10419 = ~new_n10408 & ~new_n10418;
  assign new_n10420 = ~new_n10419 & new_n5139;
  assign new_n10421 = ~new_n10398 & ~new_n10420;
  assign new_n10422 = ~new_n5011 & ~new_n10421;
  assign new_n10423 = ~new_n5207 & n3614;
  assign new_n10424 = n3646 & new_n5207;
  assign new_n10425 = ~new_n10423 & ~new_n10424;
  assign new_n10426 = ~new_n5243 & ~new_n10425;
  assign new_n10427 = ~new_n5207 & n3678;
  assign new_n10428 = n3710 & new_n5207;
  assign new_n10429 = ~new_n10427 & ~new_n10428;
  assign new_n10430 = ~new_n10429 & new_n5243;
  assign new_n10431 = ~new_n10426 & ~new_n10430;
  assign new_n10432 = ~new_n5170 & ~new_n10431;
  assign new_n10433 = ~new_n5207 & n3742;
  assign new_n10434 = n3774 & new_n5207;
  assign new_n10435 = ~new_n10433 & ~new_n10434;
  assign new_n10436 = ~new_n5243 & ~new_n10435;
  assign new_n10437 = ~new_n5207 & n3806;
  assign new_n10438 = n3838 & new_n5207;
  assign new_n10439 = ~new_n10437 & ~new_n10438;
  assign new_n10440 = ~new_n10439 & new_n5243;
  assign new_n10441 = ~new_n10436 & ~new_n10440;
  assign new_n10442 = ~new_n10441 & new_n5170;
  assign new_n10443 = ~new_n10432 & ~new_n10442;
  assign new_n10444 = ~new_n5139 & ~new_n10443;
  assign new_n10445 = ~new_n5207 & n3870;
  assign new_n10446 = n3902 & new_n5207;
  assign new_n10447 = ~new_n10445 & ~new_n10446;
  assign new_n10448 = ~new_n5243 & ~new_n10447;
  assign new_n10449 = ~new_n5207 & n3934;
  assign new_n10450 = n3966 & new_n5207;
  assign new_n10451 = ~new_n10449 & ~new_n10450;
  assign new_n10452 = ~new_n10451 & new_n5243;
  assign new_n10453 = ~new_n10448 & ~new_n10452;
  assign new_n10454 = ~new_n5170 & ~new_n10453;
  assign new_n10455 = ~new_n5207 & n3998;
  assign new_n10456 = n4030 & new_n5207;
  assign new_n10457 = ~new_n10455 & ~new_n10456;
  assign new_n10458 = ~new_n5243 & ~new_n10457;
  assign new_n10459 = ~new_n5207 & n4062;
  assign new_n10460 = n4094 & new_n5207;
  assign new_n10461 = ~new_n10459 & ~new_n10460;
  assign new_n10462 = ~new_n10461 & new_n5243;
  assign new_n10463 = ~new_n10458 & ~new_n10462;
  assign new_n10464 = ~new_n10463 & new_n5170;
  assign new_n10465 = ~new_n10454 & ~new_n10464;
  assign new_n10466 = ~new_n10465 & new_n5139;
  assign new_n10467 = ~new_n10444 & ~new_n10466;
  assign new_n10468 = ~new_n10467 & new_n5011;
  assign new_n10469 = ~new_n10422 & ~new_n10468;
  assign new_n10470 = ~new_n10469 & new_n5031;
  assign new_n10471 = ~new_n10376 & ~new_n10470;
  assign new_n10472 = ~new_n10471 & new_n5077;
  assign new_n10473 = ~new_n10282 & ~new_n10472;
  assign new_n10474 = ~new_n10473 & new_n8902;
  assign new_n10475 = ~new_n5207 & n2054;
  assign new_n10476 = n2086 & new_n5207;
  assign new_n10477 = ~new_n10475 & ~new_n10476;
  assign new_n10478 = ~new_n5243 & ~new_n10477;
  assign new_n10479 = ~new_n5207 & n2118;
  assign new_n10480 = n2150 & new_n5207;
  assign new_n10481 = ~new_n10479 & ~new_n10480;
  assign new_n10482 = ~new_n10481 & new_n5243;
  assign new_n10483 = ~new_n10478 & ~new_n10482;
  assign new_n10484 = ~new_n5170 & ~new_n10483;
  assign new_n10485 = ~new_n5207 & n2182;
  assign new_n10486 = n2214 & new_n5207;
  assign new_n10487 = ~new_n10485 & ~new_n10486;
  assign new_n10488 = ~new_n5243 & ~new_n10487;
  assign new_n10489 = ~new_n5207 & n2246;
  assign new_n10490 = n2278 & new_n5207;
  assign new_n10491 = ~new_n10489 & ~new_n10490;
  assign new_n10492 = ~new_n10491 & new_n5243;
  assign new_n10493 = ~new_n10488 & ~new_n10492;
  assign new_n10494 = ~new_n10493 & new_n5170;
  assign new_n10495 = ~new_n10484 & ~new_n10494;
  assign new_n10496 = ~new_n5139 & ~new_n10495;
  assign new_n10497 = ~new_n5207 & n2310;
  assign new_n10498 = n2342 & new_n5207;
  assign new_n10499 = ~new_n10497 & ~new_n10498;
  assign new_n10500 = ~new_n5243 & ~new_n10499;
  assign new_n10501 = ~new_n5207 & n2374;
  assign new_n10502 = n2406 & new_n5207;
  assign new_n10503 = ~new_n10501 & ~new_n10502;
  assign new_n10504 = ~new_n10503 & new_n5243;
  assign new_n10505 = ~new_n10500 & ~new_n10504;
  assign new_n10506 = ~new_n5170 & ~new_n10505;
  assign new_n10507 = ~new_n5207 & n2438;
  assign new_n10508 = n2470 & new_n5207;
  assign new_n10509 = ~new_n10507 & ~new_n10508;
  assign new_n10510 = ~new_n5243 & ~new_n10509;
  assign new_n10511 = ~new_n5207 & n2502;
  assign new_n10512 = n2534 & new_n5207;
  assign new_n10513 = ~new_n10511 & ~new_n10512;
  assign new_n10514 = ~new_n10513 & new_n5243;
  assign new_n10515 = ~new_n10510 & ~new_n10514;
  assign new_n10516 = ~new_n10515 & new_n5170;
  assign new_n10517 = ~new_n10506 & ~new_n10516;
  assign new_n10518 = ~new_n10517 & new_n5139;
  assign new_n10519 = ~new_n10496 & ~new_n10518;
  assign new_n10520 = ~new_n5011 & ~new_n10519;
  assign new_n10521 = ~new_n5207 & n2566;
  assign new_n10522 = n2598 & new_n5207;
  assign new_n10523 = ~new_n10521 & ~new_n10522;
  assign new_n10524 = ~new_n5243 & ~new_n10523;
  assign new_n10525 = ~new_n5207 & n2630;
  assign new_n10526 = n2662 & new_n5207;
  assign new_n10527 = ~new_n10525 & ~new_n10526;
  assign new_n10528 = ~new_n10527 & new_n5243;
  assign new_n10529 = ~new_n10524 & ~new_n10528;
  assign new_n10530 = ~new_n5170 & ~new_n10529;
  assign new_n10531 = ~new_n5207 & n2694;
  assign new_n10532 = n2726 & new_n5207;
  assign new_n10533 = ~new_n10531 & ~new_n10532;
  assign new_n10534 = ~new_n5243 & ~new_n10533;
  assign new_n10535 = ~new_n5207 & n2758;
  assign new_n10536 = n2790 & new_n5207;
  assign new_n10537 = ~new_n10535 & ~new_n10536;
  assign new_n10538 = ~new_n10537 & new_n5243;
  assign new_n10539 = ~new_n10534 & ~new_n10538;
  assign new_n10540 = ~new_n10539 & new_n5170;
  assign new_n10541 = ~new_n10530 & ~new_n10540;
  assign new_n10542 = ~new_n5139 & ~new_n10541;
  assign new_n10543 = ~new_n5207 & n2822;
  assign new_n10544 = n2854 & new_n5207;
  assign new_n10545 = ~new_n10543 & ~new_n10544;
  assign new_n10546 = ~new_n5243 & ~new_n10545;
  assign new_n10547 = ~new_n5207 & n2886;
  assign new_n10548 = n2918 & new_n5207;
  assign new_n10549 = ~new_n10547 & ~new_n10548;
  assign new_n10550 = ~new_n10549 & new_n5243;
  assign new_n10551 = ~new_n10546 & ~new_n10550;
  assign new_n10552 = ~new_n5170 & ~new_n10551;
  assign new_n10553 = ~new_n5207 & n2950;
  assign new_n10554 = n2982 & new_n5207;
  assign new_n10555 = ~new_n10553 & ~new_n10554;
  assign new_n10556 = ~new_n5243 & ~new_n10555;
  assign new_n10557 = ~new_n5207 & n3014;
  assign new_n10558 = n3046 & new_n5207;
  assign new_n10559 = ~new_n10557 & ~new_n10558;
  assign new_n10560 = ~new_n10559 & new_n5243;
  assign new_n10561 = ~new_n10556 & ~new_n10560;
  assign new_n10562 = ~new_n10561 & new_n5170;
  assign new_n10563 = ~new_n10552 & ~new_n10562;
  assign new_n10564 = ~new_n10563 & new_n5139;
  assign new_n10565 = ~new_n10542 & ~new_n10564;
  assign new_n10566 = ~new_n10565 & new_n5011;
  assign new_n10567 = ~new_n10520 & ~new_n10566;
  assign new_n10568 = ~new_n5031 & ~new_n10567;
  assign new_n10569 = ~new_n5207 & n3078;
  assign new_n10570 = n3110 & new_n5207;
  assign new_n10571 = ~new_n10569 & ~new_n10570;
  assign new_n10572 = ~new_n5243 & ~new_n10571;
  assign new_n10573 = ~new_n5207 & n3142;
  assign new_n10574 = n3174 & new_n5207;
  assign new_n10575 = ~new_n10573 & ~new_n10574;
  assign new_n10576 = ~new_n10575 & new_n5243;
  assign new_n10577 = ~new_n10572 & ~new_n10576;
  assign new_n10578 = ~new_n5170 & ~new_n10577;
  assign new_n10579 = ~new_n5207 & n3206;
  assign new_n10580 = n3238 & new_n5207;
  assign new_n10581 = ~new_n10579 & ~new_n10580;
  assign new_n10582 = ~new_n5243 & ~new_n10581;
  assign new_n10583 = ~new_n5207 & n3270;
  assign new_n10584 = n3302 & new_n5207;
  assign new_n10585 = ~new_n10583 & ~new_n10584;
  assign new_n10586 = ~new_n10585 & new_n5243;
  assign new_n10587 = ~new_n10582 & ~new_n10586;
  assign new_n10588 = ~new_n10587 & new_n5170;
  assign new_n10589 = ~new_n10578 & ~new_n10588;
  assign new_n10590 = ~new_n5139 & ~new_n10589;
  assign new_n10591 = ~new_n5207 & n3334;
  assign new_n10592 = n3366 & new_n5207;
  assign new_n10593 = ~new_n10591 & ~new_n10592;
  assign new_n10594 = ~new_n5243 & ~new_n10593;
  assign new_n10595 = ~new_n5207 & n3398;
  assign new_n10596 = n3430 & new_n5207;
  assign new_n10597 = ~new_n10595 & ~new_n10596;
  assign new_n10598 = ~new_n10597 & new_n5243;
  assign new_n10599 = ~new_n10594 & ~new_n10598;
  assign new_n10600 = ~new_n5170 & ~new_n10599;
  assign new_n10601 = ~new_n5207 & n3462;
  assign new_n10602 = n3494 & new_n5207;
  assign new_n10603 = ~new_n10601 & ~new_n10602;
  assign new_n10604 = ~new_n5243 & ~new_n10603;
  assign new_n10605 = ~new_n5207 & n3526;
  assign new_n10606 = n3558 & new_n5207;
  assign new_n10607 = ~new_n10605 & ~new_n10606;
  assign new_n10608 = ~new_n10607 & new_n5243;
  assign new_n10609 = ~new_n10604 & ~new_n10608;
  assign new_n10610 = ~new_n10609 & new_n5170;
  assign new_n10611 = ~new_n10600 & ~new_n10610;
  assign new_n10612 = ~new_n10611 & new_n5139;
  assign new_n10613 = ~new_n10590 & ~new_n10612;
  assign new_n10614 = ~new_n5011 & ~new_n10613;
  assign new_n10615 = ~new_n5207 & n3590;
  assign new_n10616 = n3622 & new_n5207;
  assign new_n10617 = ~new_n10615 & ~new_n10616;
  assign new_n10618 = ~new_n5243 & ~new_n10617;
  assign new_n10619 = ~new_n5207 & n3654;
  assign new_n10620 = n3686 & new_n5207;
  assign new_n10621 = ~new_n10619 & ~new_n10620;
  assign new_n10622 = ~new_n10621 & new_n5243;
  assign new_n10623 = ~new_n10618 & ~new_n10622;
  assign new_n10624 = ~new_n5170 & ~new_n10623;
  assign new_n10625 = ~new_n5207 & n3718;
  assign new_n10626 = n3750 & new_n5207;
  assign new_n10627 = ~new_n10625 & ~new_n10626;
  assign new_n10628 = ~new_n5243 & ~new_n10627;
  assign new_n10629 = ~new_n5207 & n3782;
  assign new_n10630 = n3814 & new_n5207;
  assign new_n10631 = ~new_n10629 & ~new_n10630;
  assign new_n10632 = ~new_n10631 & new_n5243;
  assign new_n10633 = ~new_n10628 & ~new_n10632;
  assign new_n10634 = ~new_n10633 & new_n5170;
  assign new_n10635 = ~new_n10624 & ~new_n10634;
  assign new_n10636 = ~new_n5139 & ~new_n10635;
  assign new_n10637 = ~new_n5207 & n3846;
  assign new_n10638 = n3878 & new_n5207;
  assign new_n10639 = ~new_n10637 & ~new_n10638;
  assign new_n10640 = ~new_n5243 & ~new_n10639;
  assign new_n10641 = ~new_n5207 & n3910;
  assign new_n10642 = n3942 & new_n5207;
  assign new_n10643 = ~new_n10641 & ~new_n10642;
  assign new_n10644 = ~new_n10643 & new_n5243;
  assign new_n10645 = ~new_n10640 & ~new_n10644;
  assign new_n10646 = ~new_n5170 & ~new_n10645;
  assign new_n10647 = ~new_n5207 & n3974;
  assign new_n10648 = n4006 & new_n5207;
  assign new_n10649 = ~new_n10647 & ~new_n10648;
  assign new_n10650 = ~new_n5243 & ~new_n10649;
  assign new_n10651 = ~new_n5207 & n4038;
  assign new_n10652 = n4070 & new_n5207;
  assign new_n10653 = ~new_n10651 & ~new_n10652;
  assign new_n10654 = ~new_n10653 & new_n5243;
  assign new_n10655 = ~new_n10650 & ~new_n10654;
  assign new_n10656 = ~new_n10655 & new_n5170;
  assign new_n10657 = ~new_n10646 & ~new_n10656;
  assign new_n10658 = ~new_n10657 & new_n5139;
  assign new_n10659 = ~new_n10636 & ~new_n10658;
  assign new_n10660 = ~new_n10659 & new_n5011;
  assign new_n10661 = ~new_n10614 & ~new_n10660;
  assign new_n10662 = ~new_n10661 & new_n5031;
  assign new_n10663 = ~new_n10568 & ~new_n10662;
  assign new_n10664 = ~new_n10663 & new_n5114;
  assign new_n10665 = ~new_n5462 & ~new_n10281;
  assign new_n10666 = ~new_n10664 & ~new_n10665;
  assign new_n10667 = ~new_n5207 & n2070;
  assign new_n10668 = n2102 & new_n5207;
  assign new_n10669 = ~new_n10667 & ~new_n10668;
  assign new_n10670 = ~new_n5243 & ~new_n10669;
  assign new_n10671 = ~new_n5207 & n2134;
  assign new_n10672 = n2166 & new_n5207;
  assign new_n10673 = ~new_n10671 & ~new_n10672;
  assign new_n10674 = ~new_n10673 & new_n5243;
  assign new_n10675 = ~new_n10670 & ~new_n10674;
  assign new_n10676 = ~new_n5170 & ~new_n10675;
  assign new_n10677 = ~new_n5207 & n2198;
  assign new_n10678 = n2230 & new_n5207;
  assign new_n10679 = ~new_n10677 & ~new_n10678;
  assign new_n10680 = ~new_n5243 & ~new_n10679;
  assign new_n10681 = ~new_n5207 & n2262;
  assign new_n10682 = n2294 & new_n5207;
  assign new_n10683 = ~new_n10681 & ~new_n10682;
  assign new_n10684 = ~new_n10683 & new_n5243;
  assign new_n10685 = ~new_n10680 & ~new_n10684;
  assign new_n10686 = ~new_n10685 & new_n5170;
  assign new_n10687 = ~new_n10676 & ~new_n10686;
  assign new_n10688 = ~new_n5139 & ~new_n10687;
  assign new_n10689 = ~new_n5207 & n2326;
  assign new_n10690 = n2358 & new_n5207;
  assign new_n10691 = ~new_n10689 & ~new_n10690;
  assign new_n10692 = ~new_n5243 & ~new_n10691;
  assign new_n10693 = ~new_n5207 & n2390;
  assign new_n10694 = n2422 & new_n5207;
  assign new_n10695 = ~new_n10693 & ~new_n10694;
  assign new_n10696 = ~new_n10695 & new_n5243;
  assign new_n10697 = ~new_n10692 & ~new_n10696;
  assign new_n10698 = ~new_n5170 & ~new_n10697;
  assign new_n10699 = ~new_n5207 & n2454;
  assign new_n10700 = n2486 & new_n5207;
  assign new_n10701 = ~new_n10699 & ~new_n10700;
  assign new_n10702 = ~new_n5243 & ~new_n10701;
  assign new_n10703 = ~new_n5207 & n2518;
  assign new_n10704 = n2550 & new_n5207;
  assign new_n10705 = ~new_n10703 & ~new_n10704;
  assign new_n10706 = ~new_n10705 & new_n5243;
  assign new_n10707 = ~new_n10702 & ~new_n10706;
  assign new_n10708 = ~new_n10707 & new_n5170;
  assign new_n10709 = ~new_n10698 & ~new_n10708;
  assign new_n10710 = ~new_n10709 & new_n5139;
  assign new_n10711 = ~new_n10688 & ~new_n10710;
  assign new_n10712 = ~new_n5011 & ~new_n10711;
  assign new_n10713 = ~new_n5207 & n2582;
  assign new_n10714 = n2614 & new_n5207;
  assign new_n10715 = ~new_n10713 & ~new_n10714;
  assign new_n10716 = ~new_n5243 & ~new_n10715;
  assign new_n10717 = ~new_n5207 & n2646;
  assign new_n10718 = n2678 & new_n5207;
  assign new_n10719 = ~new_n10717 & ~new_n10718;
  assign new_n10720 = ~new_n10719 & new_n5243;
  assign new_n10721 = ~new_n10716 & ~new_n10720;
  assign new_n10722 = ~new_n5170 & ~new_n10721;
  assign new_n10723 = ~new_n5207 & n2710;
  assign new_n10724 = n2742 & new_n5207;
  assign new_n10725 = ~new_n10723 & ~new_n10724;
  assign new_n10726 = ~new_n5243 & ~new_n10725;
  assign new_n10727 = ~new_n5207 & n2774;
  assign new_n10728 = n2806 & new_n5207;
  assign new_n10729 = ~new_n10727 & ~new_n10728;
  assign new_n10730 = ~new_n10729 & new_n5243;
  assign new_n10731 = ~new_n10726 & ~new_n10730;
  assign new_n10732 = ~new_n10731 & new_n5170;
  assign new_n10733 = ~new_n10722 & ~new_n10732;
  assign new_n10734 = ~new_n5139 & ~new_n10733;
  assign new_n10735 = ~new_n5207 & n2838;
  assign new_n10736 = n2870 & new_n5207;
  assign new_n10737 = ~new_n10735 & ~new_n10736;
  assign new_n10738 = ~new_n5243 & ~new_n10737;
  assign new_n10739 = ~new_n5207 & n2902;
  assign new_n10740 = n2934 & new_n5207;
  assign new_n10741 = ~new_n10739 & ~new_n10740;
  assign new_n10742 = ~new_n10741 & new_n5243;
  assign new_n10743 = ~new_n10738 & ~new_n10742;
  assign new_n10744 = ~new_n5170 & ~new_n10743;
  assign new_n10745 = ~new_n5207 & n2966;
  assign new_n10746 = n2998 & new_n5207;
  assign new_n10747 = ~new_n10745 & ~new_n10746;
  assign new_n10748 = ~new_n5243 & ~new_n10747;
  assign new_n10749 = ~new_n5207 & n3030;
  assign new_n10750 = n3062 & new_n5207;
  assign new_n10751 = ~new_n10749 & ~new_n10750;
  assign new_n10752 = ~new_n10751 & new_n5243;
  assign new_n10753 = ~new_n10748 & ~new_n10752;
  assign new_n10754 = ~new_n10753 & new_n5170;
  assign new_n10755 = ~new_n10744 & ~new_n10754;
  assign new_n10756 = ~new_n10755 & new_n5139;
  assign new_n10757 = ~new_n10734 & ~new_n10756;
  assign new_n10758 = ~new_n10757 & new_n5011;
  assign new_n10759 = ~new_n10712 & ~new_n10758;
  assign new_n10760 = ~new_n5031 & ~new_n10759;
  assign new_n10761 = ~new_n5207 & n3094;
  assign new_n10762 = n3126 & new_n5207;
  assign new_n10763 = ~new_n10761 & ~new_n10762;
  assign new_n10764 = ~new_n5243 & ~new_n10763;
  assign new_n10765 = ~new_n5207 & n3158;
  assign new_n10766 = n3190 & new_n5207;
  assign new_n10767 = ~new_n10765 & ~new_n10766;
  assign new_n10768 = ~new_n10767 & new_n5243;
  assign new_n10769 = ~new_n10764 & ~new_n10768;
  assign new_n10770 = ~new_n5170 & ~new_n10769;
  assign new_n10771 = ~new_n5207 & n3222;
  assign new_n10772 = n3254 & new_n5207;
  assign new_n10773 = ~new_n10771 & ~new_n10772;
  assign new_n10774 = ~new_n5243 & ~new_n10773;
  assign new_n10775 = ~new_n5207 & n3286;
  assign new_n10776 = n3318 & new_n5207;
  assign new_n10777 = ~new_n10775 & ~new_n10776;
  assign new_n10778 = ~new_n10777 & new_n5243;
  assign new_n10779 = ~new_n10774 & ~new_n10778;
  assign new_n10780 = ~new_n10779 & new_n5170;
  assign new_n10781 = ~new_n10770 & ~new_n10780;
  assign new_n10782 = ~new_n5139 & ~new_n10781;
  assign new_n10783 = ~new_n5207 & n3350;
  assign new_n10784 = n3382 & new_n5207;
  assign new_n10785 = ~new_n10783 & ~new_n10784;
  assign new_n10786 = ~new_n5243 & ~new_n10785;
  assign new_n10787 = ~new_n5207 & n3414;
  assign new_n10788 = n3446 & new_n5207;
  assign new_n10789 = ~new_n10787 & ~new_n10788;
  assign new_n10790 = ~new_n10789 & new_n5243;
  assign new_n10791 = ~new_n10786 & ~new_n10790;
  assign new_n10792 = ~new_n5170 & ~new_n10791;
  assign new_n10793 = ~new_n5207 & n3478;
  assign new_n10794 = n3510 & new_n5207;
  assign new_n10795 = ~new_n10793 & ~new_n10794;
  assign new_n10796 = ~new_n5243 & ~new_n10795;
  assign new_n10797 = ~new_n5207 & n3542;
  assign new_n10798 = n3574 & new_n5207;
  assign new_n10799 = ~new_n10797 & ~new_n10798;
  assign new_n10800 = ~new_n10799 & new_n5243;
  assign new_n10801 = ~new_n10796 & ~new_n10800;
  assign new_n10802 = ~new_n10801 & new_n5170;
  assign new_n10803 = ~new_n10792 & ~new_n10802;
  assign new_n10804 = ~new_n10803 & new_n5139;
  assign new_n10805 = ~new_n10782 & ~new_n10804;
  assign new_n10806 = ~new_n5011 & ~new_n10805;
  assign new_n10807 = ~new_n5207 & n3606;
  assign new_n10808 = n3638 & new_n5207;
  assign new_n10809 = ~new_n10807 & ~new_n10808;
  assign new_n10810 = ~new_n5243 & ~new_n10809;
  assign new_n10811 = ~new_n5207 & n3670;
  assign new_n10812 = n3702 & new_n5207;
  assign new_n10813 = ~new_n10811 & ~new_n10812;
  assign new_n10814 = ~new_n10813 & new_n5243;
  assign new_n10815 = ~new_n10810 & ~new_n10814;
  assign new_n10816 = ~new_n5170 & ~new_n10815;
  assign new_n10817 = ~new_n5207 & n3734;
  assign new_n10818 = n3766 & new_n5207;
  assign new_n10819 = ~new_n10817 & ~new_n10818;
  assign new_n10820 = ~new_n5243 & ~new_n10819;
  assign new_n10821 = ~new_n5207 & n3798;
  assign new_n10822 = n3830 & new_n5207;
  assign new_n10823 = ~new_n10821 & ~new_n10822;
  assign new_n10824 = ~new_n10823 & new_n5243;
  assign new_n10825 = ~new_n10820 & ~new_n10824;
  assign new_n10826 = ~new_n10825 & new_n5170;
  assign new_n10827 = ~new_n10816 & ~new_n10826;
  assign new_n10828 = ~new_n5139 & ~new_n10827;
  assign new_n10829 = ~new_n5207 & n3862;
  assign new_n10830 = n3894 & new_n5207;
  assign new_n10831 = ~new_n10829 & ~new_n10830;
  assign new_n10832 = ~new_n5243 & ~new_n10831;
  assign new_n10833 = ~new_n5207 & n3926;
  assign new_n10834 = n3958 & new_n5207;
  assign new_n10835 = ~new_n10833 & ~new_n10834;
  assign new_n10836 = ~new_n10835 & new_n5243;
  assign new_n10837 = ~new_n10832 & ~new_n10836;
  assign new_n10838 = ~new_n5170 & ~new_n10837;
  assign new_n10839 = ~new_n5207 & n3990;
  assign new_n10840 = n4022 & new_n5207;
  assign new_n10841 = ~new_n10839 & ~new_n10840;
  assign new_n10842 = ~new_n5243 & ~new_n10841;
  assign new_n10843 = ~new_n5207 & n4054;
  assign new_n10844 = n4086 & new_n5207;
  assign new_n10845 = ~new_n10843 & ~new_n10844;
  assign new_n10846 = ~new_n10845 & new_n5243;
  assign new_n10847 = ~new_n10842 & ~new_n10846;
  assign new_n10848 = ~new_n10847 & new_n5170;
  assign new_n10849 = ~new_n10838 & ~new_n10848;
  assign new_n10850 = ~new_n10849 & new_n5139;
  assign new_n10851 = ~new_n10828 & ~new_n10850;
  assign new_n10852 = ~new_n10851 & new_n5011;
  assign new_n10853 = ~new_n10806 & ~new_n10852;
  assign new_n10854 = ~new_n10853 & new_n5031;
  assign new_n10855 = ~new_n10760 & ~new_n10854;
  assign new_n10856 = ~new_n5115 & ~new_n10855;
  assign new_n10857 = ~new_n5116 & ~new_n10471;
  assign new_n10858 = ~new_n10856 & ~new_n10857;
  assign new_n10859 = new_n10666 & new_n10858;
  assign new_n10860 = ~new_n9289 & ~new_n10859;
  assign new_n10861 = ~new_n10474 & ~new_n10860;
  assign new_n10862 = ~new_n10092 & new_n10861;
  assign new_n10863 = ~new_n10859 & new_n8900;
  assign new_n10864 = ~new_n10473 & new_n8901;
  assign new_n10865 = ~new_n10863 & ~new_n10864;
  assign new_n10866 = ~new_n10471 & new_n4150;
  assign new_n10867 = ~new_n5207 & ~new_n9302;
  assign new_n10868 = ~new_n10866 & ~new_n10867;
  assign new_n10869 = new_n10865 & new_n10868;
  assign new_n10870 = new_n10862 & new_n10869;
  assign new_n10871 = ~new_n10870 & new_n8515;
  assign new_n10872 = ~new_n5207 & n2061;
  assign new_n10873 = n2093 & new_n5207;
  assign new_n10874 = ~new_n10872 & ~new_n10873;
  assign new_n10875 = ~new_n5243 & ~new_n10874;
  assign new_n10876 = ~new_n5207 & n2125;
  assign new_n10877 = n2157 & new_n5207;
  assign new_n10878 = ~new_n10876 & ~new_n10877;
  assign new_n10879 = ~new_n10878 & new_n5243;
  assign new_n10880 = ~new_n10875 & ~new_n10879;
  assign new_n10881 = ~new_n5170 & ~new_n10880;
  assign new_n10882 = ~new_n5207 & n2189;
  assign new_n10883 = n2221 & new_n5207;
  assign new_n10884 = ~new_n10882 & ~new_n10883;
  assign new_n10885 = ~new_n5243 & ~new_n10884;
  assign new_n10886 = ~new_n5207 & n2253;
  assign new_n10887 = n2285 & new_n5207;
  assign new_n10888 = ~new_n10886 & ~new_n10887;
  assign new_n10889 = ~new_n10888 & new_n5243;
  assign new_n10890 = ~new_n10885 & ~new_n10889;
  assign new_n10891 = ~new_n10890 & new_n5170;
  assign new_n10892 = ~new_n10881 & ~new_n10891;
  assign new_n10893 = ~new_n5139 & ~new_n10892;
  assign new_n10894 = ~new_n5207 & n2317;
  assign new_n10895 = n2349 & new_n5207;
  assign new_n10896 = ~new_n10894 & ~new_n10895;
  assign new_n10897 = ~new_n5243 & ~new_n10896;
  assign new_n10898 = ~new_n5207 & n2381;
  assign new_n10899 = n2413 & new_n5207;
  assign new_n10900 = ~new_n10898 & ~new_n10899;
  assign new_n10901 = ~new_n10900 & new_n5243;
  assign new_n10902 = ~new_n10897 & ~new_n10901;
  assign new_n10903 = ~new_n5170 & ~new_n10902;
  assign new_n10904 = ~new_n5207 & n2445;
  assign new_n10905 = n2477 & new_n5207;
  assign new_n10906 = ~new_n10904 & ~new_n10905;
  assign new_n10907 = ~new_n5243 & ~new_n10906;
  assign new_n10908 = ~new_n5207 & n2509;
  assign new_n10909 = n2541 & new_n5207;
  assign new_n10910 = ~new_n10908 & ~new_n10909;
  assign new_n10911 = ~new_n10910 & new_n5243;
  assign new_n10912 = ~new_n10907 & ~new_n10911;
  assign new_n10913 = ~new_n10912 & new_n5170;
  assign new_n10914 = ~new_n10903 & ~new_n10913;
  assign new_n10915 = ~new_n10914 & new_n5139;
  assign new_n10916 = ~new_n10893 & ~new_n10915;
  assign new_n10917 = ~new_n5011 & ~new_n10916;
  assign new_n10918 = ~new_n5207 & n2573;
  assign new_n10919 = n2605 & new_n5207;
  assign new_n10920 = ~new_n10918 & ~new_n10919;
  assign new_n10921 = ~new_n5243 & ~new_n10920;
  assign new_n10922 = ~new_n5207 & n2637;
  assign new_n10923 = n2669 & new_n5207;
  assign new_n10924 = ~new_n10922 & ~new_n10923;
  assign new_n10925 = ~new_n10924 & new_n5243;
  assign new_n10926 = ~new_n10921 & ~new_n10925;
  assign new_n10927 = ~new_n5170 & ~new_n10926;
  assign new_n10928 = ~new_n5207 & n2701;
  assign new_n10929 = n2733 & new_n5207;
  assign new_n10930 = ~new_n10928 & ~new_n10929;
  assign new_n10931 = ~new_n5243 & ~new_n10930;
  assign new_n10932 = ~new_n5207 & n2765;
  assign new_n10933 = n2797 & new_n5207;
  assign new_n10934 = ~new_n10932 & ~new_n10933;
  assign new_n10935 = ~new_n10934 & new_n5243;
  assign new_n10936 = ~new_n10931 & ~new_n10935;
  assign new_n10937 = ~new_n10936 & new_n5170;
  assign new_n10938 = ~new_n10927 & ~new_n10937;
  assign new_n10939 = ~new_n5139 & ~new_n10938;
  assign new_n10940 = ~new_n5207 & n2829;
  assign new_n10941 = n2861 & new_n5207;
  assign new_n10942 = ~new_n10940 & ~new_n10941;
  assign new_n10943 = ~new_n5243 & ~new_n10942;
  assign new_n10944 = ~new_n5207 & n2893;
  assign new_n10945 = n2925 & new_n5207;
  assign new_n10946 = ~new_n10944 & ~new_n10945;
  assign new_n10947 = ~new_n10946 & new_n5243;
  assign new_n10948 = ~new_n10943 & ~new_n10947;
  assign new_n10949 = ~new_n5170 & ~new_n10948;
  assign new_n10950 = ~new_n5207 & n2957;
  assign new_n10951 = n2989 & new_n5207;
  assign new_n10952 = ~new_n10950 & ~new_n10951;
  assign new_n10953 = ~new_n5243 & ~new_n10952;
  assign new_n10954 = ~new_n5207 & n3021;
  assign new_n10955 = n3053 & new_n5207;
  assign new_n10956 = ~new_n10954 & ~new_n10955;
  assign new_n10957 = ~new_n10956 & new_n5243;
  assign new_n10958 = ~new_n10953 & ~new_n10957;
  assign new_n10959 = ~new_n10958 & new_n5170;
  assign new_n10960 = ~new_n10949 & ~new_n10959;
  assign new_n10961 = ~new_n10960 & new_n5139;
  assign new_n10962 = ~new_n10939 & ~new_n10961;
  assign new_n10963 = ~new_n10962 & new_n5011;
  assign new_n10964 = ~new_n10917 & ~new_n10963;
  assign new_n10965 = ~new_n5031 & ~new_n10964;
  assign new_n10966 = ~new_n5207 & n3085;
  assign new_n10967 = n3117 & new_n5207;
  assign new_n10968 = ~new_n10966 & ~new_n10967;
  assign new_n10969 = ~new_n5243 & ~new_n10968;
  assign new_n10970 = ~new_n5207 & n3149;
  assign new_n10971 = n3181 & new_n5207;
  assign new_n10972 = ~new_n10970 & ~new_n10971;
  assign new_n10973 = ~new_n10972 & new_n5243;
  assign new_n10974 = ~new_n10969 & ~new_n10973;
  assign new_n10975 = ~new_n5170 & ~new_n10974;
  assign new_n10976 = ~new_n5207 & n3213;
  assign new_n10977 = n3245 & new_n5207;
  assign new_n10978 = ~new_n10976 & ~new_n10977;
  assign new_n10979 = ~new_n5243 & ~new_n10978;
  assign new_n10980 = ~new_n5207 & n3277;
  assign new_n10981 = n3309 & new_n5207;
  assign new_n10982 = ~new_n10980 & ~new_n10981;
  assign new_n10983 = ~new_n10982 & new_n5243;
  assign new_n10984 = ~new_n10979 & ~new_n10983;
  assign new_n10985 = ~new_n10984 & new_n5170;
  assign new_n10986 = ~new_n10975 & ~new_n10985;
  assign new_n10987 = ~new_n5139 & ~new_n10986;
  assign new_n10988 = ~new_n5207 & n3341;
  assign new_n10989 = n3373 & new_n5207;
  assign new_n10990 = ~new_n10988 & ~new_n10989;
  assign new_n10991 = ~new_n5243 & ~new_n10990;
  assign new_n10992 = ~new_n5207 & n3405;
  assign new_n10993 = n3437 & new_n5207;
  assign new_n10994 = ~new_n10992 & ~new_n10993;
  assign new_n10995 = ~new_n10994 & new_n5243;
  assign new_n10996 = ~new_n10991 & ~new_n10995;
  assign new_n10997 = ~new_n5170 & ~new_n10996;
  assign new_n10998 = ~new_n5207 & n3469;
  assign new_n10999 = n3501 & new_n5207;
  assign new_n11000 = ~new_n10998 & ~new_n10999;
  assign new_n11001 = ~new_n5243 & ~new_n11000;
  assign new_n11002 = ~new_n5207 & n3533;
  assign new_n11003 = n3565 & new_n5207;
  assign new_n11004 = ~new_n11002 & ~new_n11003;
  assign new_n11005 = ~new_n11004 & new_n5243;
  assign new_n11006 = ~new_n11001 & ~new_n11005;
  assign new_n11007 = ~new_n11006 & new_n5170;
  assign new_n11008 = ~new_n10997 & ~new_n11007;
  assign new_n11009 = ~new_n11008 & new_n5139;
  assign new_n11010 = ~new_n10987 & ~new_n11009;
  assign new_n11011 = ~new_n5011 & ~new_n11010;
  assign new_n11012 = ~new_n5207 & n3597;
  assign new_n11013 = n3629 & new_n5207;
  assign new_n11014 = ~new_n11012 & ~new_n11013;
  assign new_n11015 = ~new_n5243 & ~new_n11014;
  assign new_n11016 = ~new_n5207 & n3661;
  assign new_n11017 = n3693 & new_n5207;
  assign new_n11018 = ~new_n11016 & ~new_n11017;
  assign new_n11019 = ~new_n11018 & new_n5243;
  assign new_n11020 = ~new_n11015 & ~new_n11019;
  assign new_n11021 = ~new_n5170 & ~new_n11020;
  assign new_n11022 = ~new_n5207 & n3725;
  assign new_n11023 = n3757 & new_n5207;
  assign new_n11024 = ~new_n11022 & ~new_n11023;
  assign new_n11025 = ~new_n5243 & ~new_n11024;
  assign new_n11026 = ~new_n5207 & n3789;
  assign new_n11027 = n3821 & new_n5207;
  assign new_n11028 = ~new_n11026 & ~new_n11027;
  assign new_n11029 = ~new_n11028 & new_n5243;
  assign new_n11030 = ~new_n11025 & ~new_n11029;
  assign new_n11031 = ~new_n11030 & new_n5170;
  assign new_n11032 = ~new_n11021 & ~new_n11031;
  assign new_n11033 = ~new_n5139 & ~new_n11032;
  assign new_n11034 = ~new_n5207 & n3853;
  assign new_n11035 = n3885 & new_n5207;
  assign new_n11036 = ~new_n11034 & ~new_n11035;
  assign new_n11037 = ~new_n5243 & ~new_n11036;
  assign new_n11038 = ~new_n5207 & n3917;
  assign new_n11039 = n3949 & new_n5207;
  assign new_n11040 = ~new_n11038 & ~new_n11039;
  assign new_n11041 = ~new_n11040 & new_n5243;
  assign new_n11042 = ~new_n11037 & ~new_n11041;
  assign new_n11043 = ~new_n5170 & ~new_n11042;
  assign new_n11044 = ~new_n5207 & n3981;
  assign new_n11045 = n4013 & new_n5207;
  assign new_n11046 = ~new_n11044 & ~new_n11045;
  assign new_n11047 = ~new_n5243 & ~new_n11046;
  assign new_n11048 = ~new_n5207 & n4045;
  assign new_n11049 = n4077 & new_n5207;
  assign new_n11050 = ~new_n11048 & ~new_n11049;
  assign new_n11051 = ~new_n11050 & new_n5243;
  assign new_n11052 = ~new_n11047 & ~new_n11051;
  assign new_n11053 = ~new_n11052 & new_n5170;
  assign new_n11054 = ~new_n11043 & ~new_n11053;
  assign new_n11055 = ~new_n11054 & new_n5139;
  assign new_n11056 = ~new_n11033 & ~new_n11055;
  assign new_n11057 = ~new_n11056 & new_n5011;
  assign new_n11058 = ~new_n11011 & ~new_n11057;
  assign new_n11059 = ~new_n11058 & new_n5031;
  assign new_n11060 = ~new_n10965 & ~new_n11059;
  assign new_n11061 = ~new_n5077 & ~new_n11060;
  assign new_n11062 = ~new_n5207 & n2077;
  assign new_n11063 = n2109 & new_n5207;
  assign new_n11064 = ~new_n11062 & ~new_n11063;
  assign new_n11065 = ~new_n5243 & ~new_n11064;
  assign new_n11066 = ~new_n5207 & n2141;
  assign new_n11067 = n2173 & new_n5207;
  assign new_n11068 = ~new_n11066 & ~new_n11067;
  assign new_n11069 = ~new_n11068 & new_n5243;
  assign new_n11070 = ~new_n11065 & ~new_n11069;
  assign new_n11071 = ~new_n5170 & ~new_n11070;
  assign new_n11072 = ~new_n5207 & n2205;
  assign new_n11073 = n2237 & new_n5207;
  assign new_n11074 = ~new_n11072 & ~new_n11073;
  assign new_n11075 = ~new_n5243 & ~new_n11074;
  assign new_n11076 = ~new_n5207 & n2269;
  assign new_n11077 = n2301 & new_n5207;
  assign new_n11078 = ~new_n11076 & ~new_n11077;
  assign new_n11079 = ~new_n11078 & new_n5243;
  assign new_n11080 = ~new_n11075 & ~new_n11079;
  assign new_n11081 = ~new_n11080 & new_n5170;
  assign new_n11082 = ~new_n11071 & ~new_n11081;
  assign new_n11083 = ~new_n5139 & ~new_n11082;
  assign new_n11084 = ~new_n5207 & n2333;
  assign new_n11085 = n2365 & new_n5207;
  assign new_n11086 = ~new_n11084 & ~new_n11085;
  assign new_n11087 = ~new_n5243 & ~new_n11086;
  assign new_n11088 = ~new_n5207 & n2397;
  assign new_n11089 = n2429 & new_n5207;
  assign new_n11090 = ~new_n11088 & ~new_n11089;
  assign new_n11091 = ~new_n11090 & new_n5243;
  assign new_n11092 = ~new_n11087 & ~new_n11091;
  assign new_n11093 = ~new_n5170 & ~new_n11092;
  assign new_n11094 = ~new_n5207 & n2461;
  assign new_n11095 = n2493 & new_n5207;
  assign new_n11096 = ~new_n11094 & ~new_n11095;
  assign new_n11097 = ~new_n5243 & ~new_n11096;
  assign new_n11098 = ~new_n5207 & n2525;
  assign new_n11099 = n2557 & new_n5207;
  assign new_n11100 = ~new_n11098 & ~new_n11099;
  assign new_n11101 = ~new_n11100 & new_n5243;
  assign new_n11102 = ~new_n11097 & ~new_n11101;
  assign new_n11103 = ~new_n11102 & new_n5170;
  assign new_n11104 = ~new_n11093 & ~new_n11103;
  assign new_n11105 = ~new_n11104 & new_n5139;
  assign new_n11106 = ~new_n11083 & ~new_n11105;
  assign new_n11107 = ~new_n5011 & ~new_n11106;
  assign new_n11108 = ~new_n5207 & n2589;
  assign new_n11109 = n2621 & new_n5207;
  assign new_n11110 = ~new_n11108 & ~new_n11109;
  assign new_n11111 = ~new_n5243 & ~new_n11110;
  assign new_n11112 = ~new_n5207 & n2653;
  assign new_n11113 = n2685 & new_n5207;
  assign new_n11114 = ~new_n11112 & ~new_n11113;
  assign new_n11115 = ~new_n11114 & new_n5243;
  assign new_n11116 = ~new_n11111 & ~new_n11115;
  assign new_n11117 = ~new_n5170 & ~new_n11116;
  assign new_n11118 = ~new_n5207 & n2717;
  assign new_n11119 = n2749 & new_n5207;
  assign new_n11120 = ~new_n11118 & ~new_n11119;
  assign new_n11121 = ~new_n5243 & ~new_n11120;
  assign new_n11122 = ~new_n5207 & n2781;
  assign new_n11123 = n2813 & new_n5207;
  assign new_n11124 = ~new_n11122 & ~new_n11123;
  assign new_n11125 = ~new_n11124 & new_n5243;
  assign new_n11126 = ~new_n11121 & ~new_n11125;
  assign new_n11127 = ~new_n11126 & new_n5170;
  assign new_n11128 = ~new_n11117 & ~new_n11127;
  assign new_n11129 = ~new_n5139 & ~new_n11128;
  assign new_n11130 = ~new_n5207 & n2845;
  assign new_n11131 = n2877 & new_n5207;
  assign new_n11132 = ~new_n11130 & ~new_n11131;
  assign new_n11133 = ~new_n5243 & ~new_n11132;
  assign new_n11134 = ~new_n5207 & n2909;
  assign new_n11135 = n2941 & new_n5207;
  assign new_n11136 = ~new_n11134 & ~new_n11135;
  assign new_n11137 = ~new_n11136 & new_n5243;
  assign new_n11138 = ~new_n11133 & ~new_n11137;
  assign new_n11139 = ~new_n5170 & ~new_n11138;
  assign new_n11140 = ~new_n5207 & n2973;
  assign new_n11141 = n3005 & new_n5207;
  assign new_n11142 = ~new_n11140 & ~new_n11141;
  assign new_n11143 = ~new_n5243 & ~new_n11142;
  assign new_n11144 = ~new_n5207 & n3037;
  assign new_n11145 = n3069 & new_n5207;
  assign new_n11146 = ~new_n11144 & ~new_n11145;
  assign new_n11147 = ~new_n11146 & new_n5243;
  assign new_n11148 = ~new_n11143 & ~new_n11147;
  assign new_n11149 = ~new_n11148 & new_n5170;
  assign new_n11150 = ~new_n11139 & ~new_n11149;
  assign new_n11151 = ~new_n11150 & new_n5139;
  assign new_n11152 = ~new_n11129 & ~new_n11151;
  assign new_n11153 = ~new_n11152 & new_n5011;
  assign new_n11154 = ~new_n11107 & ~new_n11153;
  assign new_n11155 = ~new_n5031 & ~new_n11154;
  assign new_n11156 = ~new_n5207 & n3101;
  assign new_n11157 = n3133 & new_n5207;
  assign new_n11158 = ~new_n11156 & ~new_n11157;
  assign new_n11159 = ~new_n5243 & ~new_n11158;
  assign new_n11160 = ~new_n5207 & n3165;
  assign new_n11161 = n3197 & new_n5207;
  assign new_n11162 = ~new_n11160 & ~new_n11161;
  assign new_n11163 = ~new_n11162 & new_n5243;
  assign new_n11164 = ~new_n11159 & ~new_n11163;
  assign new_n11165 = ~new_n5170 & ~new_n11164;
  assign new_n11166 = ~new_n5207 & n3229;
  assign new_n11167 = n3261 & new_n5207;
  assign new_n11168 = ~new_n11166 & ~new_n11167;
  assign new_n11169 = ~new_n5243 & ~new_n11168;
  assign new_n11170 = ~new_n5207 & n3293;
  assign new_n11171 = n3325 & new_n5207;
  assign new_n11172 = ~new_n11170 & ~new_n11171;
  assign new_n11173 = ~new_n11172 & new_n5243;
  assign new_n11174 = ~new_n11169 & ~new_n11173;
  assign new_n11175 = ~new_n11174 & new_n5170;
  assign new_n11176 = ~new_n11165 & ~new_n11175;
  assign new_n11177 = ~new_n5139 & ~new_n11176;
  assign new_n11178 = ~new_n5207 & n3357;
  assign new_n11179 = n3389 & new_n5207;
  assign new_n11180 = ~new_n11178 & ~new_n11179;
  assign new_n11181 = ~new_n5243 & ~new_n11180;
  assign new_n11182 = ~new_n5207 & n3421;
  assign new_n11183 = n3453 & new_n5207;
  assign new_n11184 = ~new_n11182 & ~new_n11183;
  assign new_n11185 = ~new_n11184 & new_n5243;
  assign new_n11186 = ~new_n11181 & ~new_n11185;
  assign new_n11187 = ~new_n5170 & ~new_n11186;
  assign new_n11188 = ~new_n5207 & n3485;
  assign new_n11189 = n3517 & new_n5207;
  assign new_n11190 = ~new_n11188 & ~new_n11189;
  assign new_n11191 = ~new_n5243 & ~new_n11190;
  assign new_n11192 = ~new_n5207 & n3549;
  assign new_n11193 = n3581 & new_n5207;
  assign new_n11194 = ~new_n11192 & ~new_n11193;
  assign new_n11195 = ~new_n11194 & new_n5243;
  assign new_n11196 = ~new_n11191 & ~new_n11195;
  assign new_n11197 = ~new_n11196 & new_n5170;
  assign new_n11198 = ~new_n11187 & ~new_n11197;
  assign new_n11199 = ~new_n11198 & new_n5139;
  assign new_n11200 = ~new_n11177 & ~new_n11199;
  assign new_n11201 = ~new_n5011 & ~new_n11200;
  assign new_n11202 = ~new_n5207 & n3613;
  assign new_n11203 = n3645 & new_n5207;
  assign new_n11204 = ~new_n11202 & ~new_n11203;
  assign new_n11205 = ~new_n5243 & ~new_n11204;
  assign new_n11206 = ~new_n5207 & n3677;
  assign new_n11207 = n3709 & new_n5207;
  assign new_n11208 = ~new_n11206 & ~new_n11207;
  assign new_n11209 = ~new_n11208 & new_n5243;
  assign new_n11210 = ~new_n11205 & ~new_n11209;
  assign new_n11211 = ~new_n5170 & ~new_n11210;
  assign new_n11212 = ~new_n5207 & n3741;
  assign new_n11213 = n3773 & new_n5207;
  assign new_n11214 = ~new_n11212 & ~new_n11213;
  assign new_n11215 = ~new_n5243 & ~new_n11214;
  assign new_n11216 = ~new_n5207 & n3805;
  assign new_n11217 = n3837 & new_n5207;
  assign new_n11218 = ~new_n11216 & ~new_n11217;
  assign new_n11219 = ~new_n11218 & new_n5243;
  assign new_n11220 = ~new_n11215 & ~new_n11219;
  assign new_n11221 = ~new_n11220 & new_n5170;
  assign new_n11222 = ~new_n11211 & ~new_n11221;
  assign new_n11223 = ~new_n5139 & ~new_n11222;
  assign new_n11224 = ~new_n5207 & n3869;
  assign new_n11225 = n3901 & new_n5207;
  assign new_n11226 = ~new_n11224 & ~new_n11225;
  assign new_n11227 = ~new_n5243 & ~new_n11226;
  assign new_n11228 = ~new_n5207 & n3933;
  assign new_n11229 = n3965 & new_n5207;
  assign new_n11230 = ~new_n11228 & ~new_n11229;
  assign new_n11231 = ~new_n11230 & new_n5243;
  assign new_n11232 = ~new_n11227 & ~new_n11231;
  assign new_n11233 = ~new_n5170 & ~new_n11232;
  assign new_n11234 = ~new_n5207 & n3997;
  assign new_n11235 = n4029 & new_n5207;
  assign new_n11236 = ~new_n11234 & ~new_n11235;
  assign new_n11237 = ~new_n5243 & ~new_n11236;
  assign new_n11238 = ~new_n5207 & n4061;
  assign new_n11239 = n4093 & new_n5207;
  assign new_n11240 = ~new_n11238 & ~new_n11239;
  assign new_n11241 = ~new_n11240 & new_n5243;
  assign new_n11242 = ~new_n11237 & ~new_n11241;
  assign new_n11243 = ~new_n11242 & new_n5170;
  assign new_n11244 = ~new_n11233 & ~new_n11243;
  assign new_n11245 = ~new_n11244 & new_n5139;
  assign new_n11246 = ~new_n11223 & ~new_n11245;
  assign new_n11247 = ~new_n11246 & new_n5011;
  assign new_n11248 = ~new_n11201 & ~new_n11247;
  assign new_n11249 = ~new_n11248 & new_n5031;
  assign new_n11250 = ~new_n11155 & ~new_n11249;
  assign new_n11251 = ~new_n11250 & new_n5077;
  assign new_n11252 = ~new_n11061 & ~new_n11251;
  assign new_n11253 = ~new_n11252 & new_n8902;
  assign new_n11254 = ~new_n5207 & n2053;
  assign new_n11255 = n2085 & new_n5207;
  assign new_n11256 = ~new_n11254 & ~new_n11255;
  assign new_n11257 = ~new_n5243 & ~new_n11256;
  assign new_n11258 = ~new_n5207 & n2117;
  assign new_n11259 = n2149 & new_n5207;
  assign new_n11260 = ~new_n11258 & ~new_n11259;
  assign new_n11261 = ~new_n11260 & new_n5243;
  assign new_n11262 = ~new_n11257 & ~new_n11261;
  assign new_n11263 = ~new_n5170 & ~new_n11262;
  assign new_n11264 = ~new_n5207 & n2181;
  assign new_n11265 = n2213 & new_n5207;
  assign new_n11266 = ~new_n11264 & ~new_n11265;
  assign new_n11267 = ~new_n5243 & ~new_n11266;
  assign new_n11268 = ~new_n5207 & n2245;
  assign new_n11269 = n2277 & new_n5207;
  assign new_n11270 = ~new_n11268 & ~new_n11269;
  assign new_n11271 = ~new_n11270 & new_n5243;
  assign new_n11272 = ~new_n11267 & ~new_n11271;
  assign new_n11273 = ~new_n11272 & new_n5170;
  assign new_n11274 = ~new_n11263 & ~new_n11273;
  assign new_n11275 = ~new_n5139 & ~new_n11274;
  assign new_n11276 = ~new_n5207 & n2309;
  assign new_n11277 = n2341 & new_n5207;
  assign new_n11278 = ~new_n11276 & ~new_n11277;
  assign new_n11279 = ~new_n5243 & ~new_n11278;
  assign new_n11280 = ~new_n5207 & n2373;
  assign new_n11281 = n2405 & new_n5207;
  assign new_n11282 = ~new_n11280 & ~new_n11281;
  assign new_n11283 = ~new_n11282 & new_n5243;
  assign new_n11284 = ~new_n11279 & ~new_n11283;
  assign new_n11285 = ~new_n5170 & ~new_n11284;
  assign new_n11286 = ~new_n5207 & n2437;
  assign new_n11287 = n2469 & new_n5207;
  assign new_n11288 = ~new_n11286 & ~new_n11287;
  assign new_n11289 = ~new_n5243 & ~new_n11288;
  assign new_n11290 = ~new_n5207 & n2501;
  assign new_n11291 = n2533 & new_n5207;
  assign new_n11292 = ~new_n11290 & ~new_n11291;
  assign new_n11293 = ~new_n11292 & new_n5243;
  assign new_n11294 = ~new_n11289 & ~new_n11293;
  assign new_n11295 = ~new_n11294 & new_n5170;
  assign new_n11296 = ~new_n11285 & ~new_n11295;
  assign new_n11297 = ~new_n11296 & new_n5139;
  assign new_n11298 = ~new_n11275 & ~new_n11297;
  assign new_n11299 = ~new_n5011 & ~new_n11298;
  assign new_n11300 = ~new_n5207 & n2565;
  assign new_n11301 = n2597 & new_n5207;
  assign new_n11302 = ~new_n11300 & ~new_n11301;
  assign new_n11303 = ~new_n5243 & ~new_n11302;
  assign new_n11304 = ~new_n5207 & n2629;
  assign new_n11305 = n2661 & new_n5207;
  assign new_n11306 = ~new_n11304 & ~new_n11305;
  assign new_n11307 = ~new_n11306 & new_n5243;
  assign new_n11308 = ~new_n11303 & ~new_n11307;
  assign new_n11309 = ~new_n5170 & ~new_n11308;
  assign new_n11310 = ~new_n5207 & n2693;
  assign new_n11311 = n2725 & new_n5207;
  assign new_n11312 = ~new_n11310 & ~new_n11311;
  assign new_n11313 = ~new_n5243 & ~new_n11312;
  assign new_n11314 = ~new_n5207 & n2757;
  assign new_n11315 = n2789 & new_n5207;
  assign new_n11316 = ~new_n11314 & ~new_n11315;
  assign new_n11317 = ~new_n11316 & new_n5243;
  assign new_n11318 = ~new_n11313 & ~new_n11317;
  assign new_n11319 = ~new_n11318 & new_n5170;
  assign new_n11320 = ~new_n11309 & ~new_n11319;
  assign new_n11321 = ~new_n5139 & ~new_n11320;
  assign new_n11322 = ~new_n5207 & n2821;
  assign new_n11323 = n2853 & new_n5207;
  assign new_n11324 = ~new_n11322 & ~new_n11323;
  assign new_n11325 = ~new_n5243 & ~new_n11324;
  assign new_n11326 = ~new_n5207 & n2885;
  assign new_n11327 = n2917 & new_n5207;
  assign new_n11328 = ~new_n11326 & ~new_n11327;
  assign new_n11329 = ~new_n11328 & new_n5243;
  assign new_n11330 = ~new_n11325 & ~new_n11329;
  assign new_n11331 = ~new_n5170 & ~new_n11330;
  assign new_n11332 = ~new_n5207 & n2949;
  assign new_n11333 = n2981 & new_n5207;
  assign new_n11334 = ~new_n11332 & ~new_n11333;
  assign new_n11335 = ~new_n5243 & ~new_n11334;
  assign new_n11336 = ~new_n5207 & n3013;
  assign new_n11337 = n3045 & new_n5207;
  assign new_n11338 = ~new_n11336 & ~new_n11337;
  assign new_n11339 = ~new_n11338 & new_n5243;
  assign new_n11340 = ~new_n11335 & ~new_n11339;
  assign new_n11341 = ~new_n11340 & new_n5170;
  assign new_n11342 = ~new_n11331 & ~new_n11341;
  assign new_n11343 = ~new_n11342 & new_n5139;
  assign new_n11344 = ~new_n11321 & ~new_n11343;
  assign new_n11345 = ~new_n11344 & new_n5011;
  assign new_n11346 = ~new_n11299 & ~new_n11345;
  assign new_n11347 = ~new_n5031 & ~new_n11346;
  assign new_n11348 = ~new_n5207 & n3077;
  assign new_n11349 = n3109 & new_n5207;
  assign new_n11350 = ~new_n11348 & ~new_n11349;
  assign new_n11351 = ~new_n5243 & ~new_n11350;
  assign new_n11352 = ~new_n5207 & n3141;
  assign new_n11353 = n3173 & new_n5207;
  assign new_n11354 = ~new_n11352 & ~new_n11353;
  assign new_n11355 = ~new_n11354 & new_n5243;
  assign new_n11356 = ~new_n11351 & ~new_n11355;
  assign new_n11357 = ~new_n5170 & ~new_n11356;
  assign new_n11358 = ~new_n5207 & n3205;
  assign new_n11359 = n3237 & new_n5207;
  assign new_n11360 = ~new_n11358 & ~new_n11359;
  assign new_n11361 = ~new_n5243 & ~new_n11360;
  assign new_n11362 = ~new_n5207 & n3269;
  assign new_n11363 = n3301 & new_n5207;
  assign new_n11364 = ~new_n11362 & ~new_n11363;
  assign new_n11365 = ~new_n11364 & new_n5243;
  assign new_n11366 = ~new_n11361 & ~new_n11365;
  assign new_n11367 = ~new_n11366 & new_n5170;
  assign new_n11368 = ~new_n11357 & ~new_n11367;
  assign new_n11369 = ~new_n5139 & ~new_n11368;
  assign new_n11370 = ~new_n5207 & n3333;
  assign new_n11371 = n3365 & new_n5207;
  assign new_n11372 = ~new_n11370 & ~new_n11371;
  assign new_n11373 = ~new_n5243 & ~new_n11372;
  assign new_n11374 = ~new_n5207 & n3397;
  assign new_n11375 = n3429 & new_n5207;
  assign new_n11376 = ~new_n11374 & ~new_n11375;
  assign new_n11377 = ~new_n11376 & new_n5243;
  assign new_n11378 = ~new_n11373 & ~new_n11377;
  assign new_n11379 = ~new_n5170 & ~new_n11378;
  assign new_n11380 = ~new_n5207 & n3461;
  assign new_n11381 = n3493 & new_n5207;
  assign new_n11382 = ~new_n11380 & ~new_n11381;
  assign new_n11383 = ~new_n5243 & ~new_n11382;
  assign new_n11384 = ~new_n5207 & n3525;
  assign new_n11385 = n3557 & new_n5207;
  assign new_n11386 = ~new_n11384 & ~new_n11385;
  assign new_n11387 = ~new_n11386 & new_n5243;
  assign new_n11388 = ~new_n11383 & ~new_n11387;
  assign new_n11389 = ~new_n11388 & new_n5170;
  assign new_n11390 = ~new_n11379 & ~new_n11389;
  assign new_n11391 = ~new_n11390 & new_n5139;
  assign new_n11392 = ~new_n11369 & ~new_n11391;
  assign new_n11393 = ~new_n5011 & ~new_n11392;
  assign new_n11394 = ~new_n5207 & n3589;
  assign new_n11395 = n3621 & new_n5207;
  assign new_n11396 = ~new_n11394 & ~new_n11395;
  assign new_n11397 = ~new_n5243 & ~new_n11396;
  assign new_n11398 = ~new_n5207 & n3653;
  assign new_n11399 = n3685 & new_n5207;
  assign new_n11400 = ~new_n11398 & ~new_n11399;
  assign new_n11401 = ~new_n11400 & new_n5243;
  assign new_n11402 = ~new_n11397 & ~new_n11401;
  assign new_n11403 = ~new_n5170 & ~new_n11402;
  assign new_n11404 = ~new_n5207 & n3717;
  assign new_n11405 = n3749 & new_n5207;
  assign new_n11406 = ~new_n11404 & ~new_n11405;
  assign new_n11407 = ~new_n5243 & ~new_n11406;
  assign new_n11408 = ~new_n5207 & n3781;
  assign new_n11409 = n3813 & new_n5207;
  assign new_n11410 = ~new_n11408 & ~new_n11409;
  assign new_n11411 = ~new_n11410 & new_n5243;
  assign new_n11412 = ~new_n11407 & ~new_n11411;
  assign new_n11413 = ~new_n11412 & new_n5170;
  assign new_n11414 = ~new_n11403 & ~new_n11413;
  assign new_n11415 = ~new_n5139 & ~new_n11414;
  assign new_n11416 = ~new_n5207 & n3845;
  assign new_n11417 = n3877 & new_n5207;
  assign new_n11418 = ~new_n11416 & ~new_n11417;
  assign new_n11419 = ~new_n5243 & ~new_n11418;
  assign new_n11420 = ~new_n5207 & n3909;
  assign new_n11421 = n3941 & new_n5207;
  assign new_n11422 = ~new_n11420 & ~new_n11421;
  assign new_n11423 = ~new_n11422 & new_n5243;
  assign new_n11424 = ~new_n11419 & ~new_n11423;
  assign new_n11425 = ~new_n5170 & ~new_n11424;
  assign new_n11426 = ~new_n5207 & n3973;
  assign new_n11427 = n4005 & new_n5207;
  assign new_n11428 = ~new_n11426 & ~new_n11427;
  assign new_n11429 = ~new_n5243 & ~new_n11428;
  assign new_n11430 = ~new_n5207 & n4037;
  assign new_n11431 = n4069 & new_n5207;
  assign new_n11432 = ~new_n11430 & ~new_n11431;
  assign new_n11433 = ~new_n11432 & new_n5243;
  assign new_n11434 = ~new_n11429 & ~new_n11433;
  assign new_n11435 = ~new_n11434 & new_n5170;
  assign new_n11436 = ~new_n11425 & ~new_n11435;
  assign new_n11437 = ~new_n11436 & new_n5139;
  assign new_n11438 = ~new_n11415 & ~new_n11437;
  assign new_n11439 = ~new_n11438 & new_n5011;
  assign new_n11440 = ~new_n11393 & ~new_n11439;
  assign new_n11441 = ~new_n11440 & new_n5031;
  assign new_n11442 = ~new_n11347 & ~new_n11441;
  assign new_n11443 = ~new_n11442 & new_n5114;
  assign new_n11444 = ~new_n5462 & ~new_n11060;
  assign new_n11445 = ~new_n11443 & ~new_n11444;
  assign new_n11446 = ~new_n5207 & n2069;
  assign new_n11447 = n2101 & new_n5207;
  assign new_n11448 = ~new_n11446 & ~new_n11447;
  assign new_n11449 = ~new_n5243 & ~new_n11448;
  assign new_n11450 = ~new_n5207 & n2133;
  assign new_n11451 = n2165 & new_n5207;
  assign new_n11452 = ~new_n11450 & ~new_n11451;
  assign new_n11453 = ~new_n11452 & new_n5243;
  assign new_n11454 = ~new_n11449 & ~new_n11453;
  assign new_n11455 = ~new_n5170 & ~new_n11454;
  assign new_n11456 = ~new_n5207 & n2197;
  assign new_n11457 = n2229 & new_n5207;
  assign new_n11458 = ~new_n11456 & ~new_n11457;
  assign new_n11459 = ~new_n5243 & ~new_n11458;
  assign new_n11460 = ~new_n5207 & n2261;
  assign new_n11461 = n2293 & new_n5207;
  assign new_n11462 = ~new_n11460 & ~new_n11461;
  assign new_n11463 = ~new_n11462 & new_n5243;
  assign new_n11464 = ~new_n11459 & ~new_n11463;
  assign new_n11465 = ~new_n11464 & new_n5170;
  assign new_n11466 = ~new_n11455 & ~new_n11465;
  assign new_n11467 = ~new_n5139 & ~new_n11466;
  assign new_n11468 = ~new_n5207 & n2325;
  assign new_n11469 = n2357 & new_n5207;
  assign new_n11470 = ~new_n11468 & ~new_n11469;
  assign new_n11471 = ~new_n5243 & ~new_n11470;
  assign new_n11472 = ~new_n5207 & n2389;
  assign new_n11473 = n2421 & new_n5207;
  assign new_n11474 = ~new_n11472 & ~new_n11473;
  assign new_n11475 = ~new_n11474 & new_n5243;
  assign new_n11476 = ~new_n11471 & ~new_n11475;
  assign new_n11477 = ~new_n5170 & ~new_n11476;
  assign new_n11478 = ~new_n5207 & n2453;
  assign new_n11479 = n2485 & new_n5207;
  assign new_n11480 = ~new_n11478 & ~new_n11479;
  assign new_n11481 = ~new_n5243 & ~new_n11480;
  assign new_n11482 = ~new_n5207 & n2517;
  assign new_n11483 = n2549 & new_n5207;
  assign new_n11484 = ~new_n11482 & ~new_n11483;
  assign new_n11485 = ~new_n11484 & new_n5243;
  assign new_n11486 = ~new_n11481 & ~new_n11485;
  assign new_n11487 = ~new_n11486 & new_n5170;
  assign new_n11488 = ~new_n11477 & ~new_n11487;
  assign new_n11489 = ~new_n11488 & new_n5139;
  assign new_n11490 = ~new_n11467 & ~new_n11489;
  assign new_n11491 = ~new_n5011 & ~new_n11490;
  assign new_n11492 = ~new_n5207 & n2581;
  assign new_n11493 = n2613 & new_n5207;
  assign new_n11494 = ~new_n11492 & ~new_n11493;
  assign new_n11495 = ~new_n5243 & ~new_n11494;
  assign new_n11496 = ~new_n5207 & n2645;
  assign new_n11497 = n2677 & new_n5207;
  assign new_n11498 = ~new_n11496 & ~new_n11497;
  assign new_n11499 = ~new_n11498 & new_n5243;
  assign new_n11500 = ~new_n11495 & ~new_n11499;
  assign new_n11501 = ~new_n5170 & ~new_n11500;
  assign new_n11502 = ~new_n5207 & n2709;
  assign new_n11503 = n2741 & new_n5207;
  assign new_n11504 = ~new_n11502 & ~new_n11503;
  assign new_n11505 = ~new_n5243 & ~new_n11504;
  assign new_n11506 = ~new_n5207 & n2773;
  assign new_n11507 = n2805 & new_n5207;
  assign new_n11508 = ~new_n11506 & ~new_n11507;
  assign new_n11509 = ~new_n11508 & new_n5243;
  assign new_n11510 = ~new_n11505 & ~new_n11509;
  assign new_n11511 = ~new_n11510 & new_n5170;
  assign new_n11512 = ~new_n11501 & ~new_n11511;
  assign new_n11513 = ~new_n5139 & ~new_n11512;
  assign new_n11514 = ~new_n5207 & n2837;
  assign new_n11515 = n2869 & new_n5207;
  assign new_n11516 = ~new_n11514 & ~new_n11515;
  assign new_n11517 = ~new_n5243 & ~new_n11516;
  assign new_n11518 = ~new_n5207 & n2901;
  assign new_n11519 = n2933 & new_n5207;
  assign new_n11520 = ~new_n11518 & ~new_n11519;
  assign new_n11521 = ~new_n11520 & new_n5243;
  assign new_n11522 = ~new_n11517 & ~new_n11521;
  assign new_n11523 = ~new_n5170 & ~new_n11522;
  assign new_n11524 = ~new_n5207 & n2965;
  assign new_n11525 = n2997 & new_n5207;
  assign new_n11526 = ~new_n11524 & ~new_n11525;
  assign new_n11527 = ~new_n5243 & ~new_n11526;
  assign new_n11528 = ~new_n5207 & n3029;
  assign new_n11529 = n3061 & new_n5207;
  assign new_n11530 = ~new_n11528 & ~new_n11529;
  assign new_n11531 = ~new_n11530 & new_n5243;
  assign new_n11532 = ~new_n11527 & ~new_n11531;
  assign new_n11533 = ~new_n11532 & new_n5170;
  assign new_n11534 = ~new_n11523 & ~new_n11533;
  assign new_n11535 = ~new_n11534 & new_n5139;
  assign new_n11536 = ~new_n11513 & ~new_n11535;
  assign new_n11537 = ~new_n11536 & new_n5011;
  assign new_n11538 = ~new_n11491 & ~new_n11537;
  assign new_n11539 = ~new_n5031 & ~new_n11538;
  assign new_n11540 = ~new_n5207 & n3093;
  assign new_n11541 = n3125 & new_n5207;
  assign new_n11542 = ~new_n11540 & ~new_n11541;
  assign new_n11543 = ~new_n5243 & ~new_n11542;
  assign new_n11544 = ~new_n5207 & n3157;
  assign new_n11545 = n3189 & new_n5207;
  assign new_n11546 = ~new_n11544 & ~new_n11545;
  assign new_n11547 = ~new_n11546 & new_n5243;
  assign new_n11548 = ~new_n11543 & ~new_n11547;
  assign new_n11549 = ~new_n5170 & ~new_n11548;
  assign new_n11550 = ~new_n5207 & n3221;
  assign new_n11551 = n3253 & new_n5207;
  assign new_n11552 = ~new_n11550 & ~new_n11551;
  assign new_n11553 = ~new_n5243 & ~new_n11552;
  assign new_n11554 = ~new_n5207 & n3285;
  assign new_n11555 = n3317 & new_n5207;
  assign new_n11556 = ~new_n11554 & ~new_n11555;
  assign new_n11557 = ~new_n11556 & new_n5243;
  assign new_n11558 = ~new_n11553 & ~new_n11557;
  assign new_n11559 = ~new_n11558 & new_n5170;
  assign new_n11560 = ~new_n11549 & ~new_n11559;
  assign new_n11561 = ~new_n5139 & ~new_n11560;
  assign new_n11562 = ~new_n5207 & n3349;
  assign new_n11563 = n3381 & new_n5207;
  assign new_n11564 = ~new_n11562 & ~new_n11563;
  assign new_n11565 = ~new_n5243 & ~new_n11564;
  assign new_n11566 = ~new_n5207 & n3413;
  assign new_n11567 = n3445 & new_n5207;
  assign new_n11568 = ~new_n11566 & ~new_n11567;
  assign new_n11569 = ~new_n11568 & new_n5243;
  assign new_n11570 = ~new_n11565 & ~new_n11569;
  assign new_n11571 = ~new_n5170 & ~new_n11570;
  assign new_n11572 = ~new_n5207 & n3477;
  assign new_n11573 = n3509 & new_n5207;
  assign new_n11574 = ~new_n11572 & ~new_n11573;
  assign new_n11575 = ~new_n5243 & ~new_n11574;
  assign new_n11576 = ~new_n5207 & n3541;
  assign new_n11577 = n3573 & new_n5207;
  assign new_n11578 = ~new_n11576 & ~new_n11577;
  assign new_n11579 = ~new_n11578 & new_n5243;
  assign new_n11580 = ~new_n11575 & ~new_n11579;
  assign new_n11581 = ~new_n11580 & new_n5170;
  assign new_n11582 = ~new_n11571 & ~new_n11581;
  assign new_n11583 = ~new_n11582 & new_n5139;
  assign new_n11584 = ~new_n11561 & ~new_n11583;
  assign new_n11585 = ~new_n5011 & ~new_n11584;
  assign new_n11586 = ~new_n5207 & n3605;
  assign new_n11587 = n3637 & new_n5207;
  assign new_n11588 = ~new_n11586 & ~new_n11587;
  assign new_n11589 = ~new_n5243 & ~new_n11588;
  assign new_n11590 = ~new_n5207 & n3669;
  assign new_n11591 = n3701 & new_n5207;
  assign new_n11592 = ~new_n11590 & ~new_n11591;
  assign new_n11593 = ~new_n11592 & new_n5243;
  assign new_n11594 = ~new_n11589 & ~new_n11593;
  assign new_n11595 = ~new_n5170 & ~new_n11594;
  assign new_n11596 = ~new_n5207 & n3733;
  assign new_n11597 = n3765 & new_n5207;
  assign new_n11598 = ~new_n11596 & ~new_n11597;
  assign new_n11599 = ~new_n5243 & ~new_n11598;
  assign new_n11600 = ~new_n5207 & n3797;
  assign new_n11601 = n3829 & new_n5207;
  assign new_n11602 = ~new_n11600 & ~new_n11601;
  assign new_n11603 = ~new_n11602 & new_n5243;
  assign new_n11604 = ~new_n11599 & ~new_n11603;
  assign new_n11605 = ~new_n11604 & new_n5170;
  assign new_n11606 = ~new_n11595 & ~new_n11605;
  assign new_n11607 = ~new_n5139 & ~new_n11606;
  assign new_n11608 = ~new_n5207 & n3861;
  assign new_n11609 = n3893 & new_n5207;
  assign new_n11610 = ~new_n11608 & ~new_n11609;
  assign new_n11611 = ~new_n5243 & ~new_n11610;
  assign new_n11612 = ~new_n5207 & n3925;
  assign new_n11613 = n3957 & new_n5207;
  assign new_n11614 = ~new_n11612 & ~new_n11613;
  assign new_n11615 = ~new_n11614 & new_n5243;
  assign new_n11616 = ~new_n11611 & ~new_n11615;
  assign new_n11617 = ~new_n5170 & ~new_n11616;
  assign new_n11618 = ~new_n5207 & n3989;
  assign new_n11619 = n4021 & new_n5207;
  assign new_n11620 = ~new_n11618 & ~new_n11619;
  assign new_n11621 = ~new_n5243 & ~new_n11620;
  assign new_n11622 = ~new_n5207 & n4053;
  assign new_n11623 = n4085 & new_n5207;
  assign new_n11624 = ~new_n11622 & ~new_n11623;
  assign new_n11625 = ~new_n11624 & new_n5243;
  assign new_n11626 = ~new_n11621 & ~new_n11625;
  assign new_n11627 = ~new_n11626 & new_n5170;
  assign new_n11628 = ~new_n11617 & ~new_n11627;
  assign new_n11629 = ~new_n11628 & new_n5139;
  assign new_n11630 = ~new_n11607 & ~new_n11629;
  assign new_n11631 = ~new_n11630 & new_n5011;
  assign new_n11632 = ~new_n11585 & ~new_n11631;
  assign new_n11633 = ~new_n11632 & new_n5031;
  assign new_n11634 = ~new_n11539 & ~new_n11633;
  assign new_n11635 = ~new_n5115 & ~new_n11634;
  assign new_n11636 = ~new_n5116 & ~new_n11250;
  assign new_n11637 = ~new_n11635 & ~new_n11636;
  assign new_n11638 = new_n11445 & new_n11637;
  assign new_n11639 = ~new_n9289 & ~new_n11638;
  assign new_n11640 = ~new_n11253 & ~new_n11639;
  assign new_n11641 = ~new_n11638 & new_n8900;
  assign new_n11642 = ~new_n11252 & new_n8901;
  assign new_n11643 = ~new_n11641 & ~new_n11642;
  assign new_n11644 = ~new_n11250 & new_n4150;
  assign new_n11645 = ~new_n5243 & ~new_n9302;
  assign new_n11646 = ~new_n11644 & ~new_n11645;
  assign new_n11647 = new_n11643 & new_n11646;
  assign new_n11648 = new_n11640 & new_n11647;
  assign new_n11649 = ~new_n11648 & new_n8515;
  assign new_n11650 = ~new_n5207 & n2060;
  assign new_n11651 = n2092 & new_n5207;
  assign new_n11652 = ~new_n11650 & ~new_n11651;
  assign new_n11653 = ~new_n5243 & ~new_n11652;
  assign new_n11654 = ~new_n5207 & n2124;
  assign new_n11655 = n2156 & new_n5207;
  assign new_n11656 = ~new_n11654 & ~new_n11655;
  assign new_n11657 = ~new_n11656 & new_n5243;
  assign new_n11658 = ~new_n11653 & ~new_n11657;
  assign new_n11659 = ~new_n5170 & ~new_n11658;
  assign new_n11660 = ~new_n5207 & n2188;
  assign new_n11661 = n2220 & new_n5207;
  assign new_n11662 = ~new_n11660 & ~new_n11661;
  assign new_n11663 = ~new_n5243 & ~new_n11662;
  assign new_n11664 = ~new_n5207 & n2252;
  assign new_n11665 = n2284 & new_n5207;
  assign new_n11666 = ~new_n11664 & ~new_n11665;
  assign new_n11667 = ~new_n11666 & new_n5243;
  assign new_n11668 = ~new_n11663 & ~new_n11667;
  assign new_n11669 = ~new_n11668 & new_n5170;
  assign new_n11670 = ~new_n11659 & ~new_n11669;
  assign new_n11671 = ~new_n5139 & ~new_n11670;
  assign new_n11672 = ~new_n5207 & n2316;
  assign new_n11673 = n2348 & new_n5207;
  assign new_n11674 = ~new_n11672 & ~new_n11673;
  assign new_n11675 = ~new_n5243 & ~new_n11674;
  assign new_n11676 = ~new_n5207 & n2380;
  assign new_n11677 = n2412 & new_n5207;
  assign new_n11678 = ~new_n11676 & ~new_n11677;
  assign new_n11679 = ~new_n11678 & new_n5243;
  assign new_n11680 = ~new_n11675 & ~new_n11679;
  assign new_n11681 = ~new_n5170 & ~new_n11680;
  assign new_n11682 = ~new_n5207 & n2444;
  assign new_n11683 = n2476 & new_n5207;
  assign new_n11684 = ~new_n11682 & ~new_n11683;
  assign new_n11685 = ~new_n5243 & ~new_n11684;
  assign new_n11686 = ~new_n5207 & n2508;
  assign new_n11687 = n2540 & new_n5207;
  assign new_n11688 = ~new_n11686 & ~new_n11687;
  assign new_n11689 = ~new_n11688 & new_n5243;
  assign new_n11690 = ~new_n11685 & ~new_n11689;
  assign new_n11691 = ~new_n11690 & new_n5170;
  assign new_n11692 = ~new_n11681 & ~new_n11691;
  assign new_n11693 = ~new_n11692 & new_n5139;
  assign new_n11694 = ~new_n11671 & ~new_n11693;
  assign new_n11695 = ~new_n5011 & ~new_n11694;
  assign new_n11696 = ~new_n5207 & n2572;
  assign new_n11697 = n2604 & new_n5207;
  assign new_n11698 = ~new_n11696 & ~new_n11697;
  assign new_n11699 = ~new_n5243 & ~new_n11698;
  assign new_n11700 = ~new_n5207 & n2636;
  assign new_n11701 = n2668 & new_n5207;
  assign new_n11702 = ~new_n11700 & ~new_n11701;
  assign new_n11703 = ~new_n11702 & new_n5243;
  assign new_n11704 = ~new_n11699 & ~new_n11703;
  assign new_n11705 = ~new_n5170 & ~new_n11704;
  assign new_n11706 = ~new_n5207 & n2700;
  assign new_n11707 = n2732 & new_n5207;
  assign new_n11708 = ~new_n11706 & ~new_n11707;
  assign new_n11709 = ~new_n5243 & ~new_n11708;
  assign new_n11710 = ~new_n5207 & n2764;
  assign new_n11711 = n2796 & new_n5207;
  assign new_n11712 = ~new_n11710 & ~new_n11711;
  assign new_n11713 = ~new_n11712 & new_n5243;
  assign new_n11714 = ~new_n11709 & ~new_n11713;
  assign new_n11715 = ~new_n11714 & new_n5170;
  assign new_n11716 = ~new_n11705 & ~new_n11715;
  assign new_n11717 = ~new_n5139 & ~new_n11716;
  assign new_n11718 = ~new_n5207 & n2828;
  assign new_n11719 = n2860 & new_n5207;
  assign new_n11720 = ~new_n11718 & ~new_n11719;
  assign new_n11721 = ~new_n5243 & ~new_n11720;
  assign new_n11722 = ~new_n5207 & n2892;
  assign new_n11723 = n2924 & new_n5207;
  assign new_n11724 = ~new_n11722 & ~new_n11723;
  assign new_n11725 = ~new_n11724 & new_n5243;
  assign new_n11726 = ~new_n11721 & ~new_n11725;
  assign new_n11727 = ~new_n5170 & ~new_n11726;
  assign new_n11728 = ~new_n5207 & n2956;
  assign new_n11729 = n2988 & new_n5207;
  assign new_n11730 = ~new_n11728 & ~new_n11729;
  assign new_n11731 = ~new_n5243 & ~new_n11730;
  assign new_n11732 = ~new_n5207 & n3020;
  assign new_n11733 = n3052 & new_n5207;
  assign new_n11734 = ~new_n11732 & ~new_n11733;
  assign new_n11735 = ~new_n11734 & new_n5243;
  assign new_n11736 = ~new_n11731 & ~new_n11735;
  assign new_n11737 = ~new_n11736 & new_n5170;
  assign new_n11738 = ~new_n11727 & ~new_n11737;
  assign new_n11739 = ~new_n11738 & new_n5139;
  assign new_n11740 = ~new_n11717 & ~new_n11739;
  assign new_n11741 = ~new_n11740 & new_n5011;
  assign new_n11742 = ~new_n11695 & ~new_n11741;
  assign new_n11743 = ~new_n5031 & ~new_n11742;
  assign new_n11744 = ~new_n5207 & n3084;
  assign new_n11745 = n3116 & new_n5207;
  assign new_n11746 = ~new_n11744 & ~new_n11745;
  assign new_n11747 = ~new_n5243 & ~new_n11746;
  assign new_n11748 = ~new_n5207 & n3148;
  assign new_n11749 = n3180 & new_n5207;
  assign new_n11750 = ~new_n11748 & ~new_n11749;
  assign new_n11751 = ~new_n11750 & new_n5243;
  assign new_n11752 = ~new_n11747 & ~new_n11751;
  assign new_n11753 = ~new_n5170 & ~new_n11752;
  assign new_n11754 = ~new_n5207 & n3212;
  assign new_n11755 = n3244 & new_n5207;
  assign new_n11756 = ~new_n11754 & ~new_n11755;
  assign new_n11757 = ~new_n5243 & ~new_n11756;
  assign new_n11758 = ~new_n5207 & n3276;
  assign new_n11759 = n3308 & new_n5207;
  assign new_n11760 = ~new_n11758 & ~new_n11759;
  assign new_n11761 = ~new_n11760 & new_n5243;
  assign new_n11762 = ~new_n11757 & ~new_n11761;
  assign new_n11763 = ~new_n11762 & new_n5170;
  assign new_n11764 = ~new_n11753 & ~new_n11763;
  assign new_n11765 = ~new_n5139 & ~new_n11764;
  assign new_n11766 = ~new_n5207 & n3340;
  assign new_n11767 = n3372 & new_n5207;
  assign new_n11768 = ~new_n11766 & ~new_n11767;
  assign new_n11769 = ~new_n5243 & ~new_n11768;
  assign new_n11770 = ~new_n5207 & n3404;
  assign new_n11771 = n3436 & new_n5207;
  assign new_n11772 = ~new_n11770 & ~new_n11771;
  assign new_n11773 = ~new_n11772 & new_n5243;
  assign new_n11774 = ~new_n11769 & ~new_n11773;
  assign new_n11775 = ~new_n5170 & ~new_n11774;
  assign new_n11776 = ~new_n5207 & n3468;
  assign new_n11777 = n3500 & new_n5207;
  assign new_n11778 = ~new_n11776 & ~new_n11777;
  assign new_n11779 = ~new_n5243 & ~new_n11778;
  assign new_n11780 = ~new_n5207 & n3532;
  assign new_n11781 = n3564 & new_n5207;
  assign new_n11782 = ~new_n11780 & ~new_n11781;
  assign new_n11783 = ~new_n11782 & new_n5243;
  assign new_n11784 = ~new_n11779 & ~new_n11783;
  assign new_n11785 = ~new_n11784 & new_n5170;
  assign new_n11786 = ~new_n11775 & ~new_n11785;
  assign new_n11787 = ~new_n11786 & new_n5139;
  assign new_n11788 = ~new_n11765 & ~new_n11787;
  assign new_n11789 = ~new_n5011 & ~new_n11788;
  assign new_n11790 = ~new_n5207 & n3596;
  assign new_n11791 = n3628 & new_n5207;
  assign new_n11792 = ~new_n11790 & ~new_n11791;
  assign new_n11793 = ~new_n5243 & ~new_n11792;
  assign new_n11794 = ~new_n5207 & n3660;
  assign new_n11795 = n3692 & new_n5207;
  assign new_n11796 = ~new_n11794 & ~new_n11795;
  assign new_n11797 = ~new_n11796 & new_n5243;
  assign new_n11798 = ~new_n11793 & ~new_n11797;
  assign new_n11799 = ~new_n5170 & ~new_n11798;
  assign new_n11800 = ~new_n5207 & n3724;
  assign new_n11801 = n3756 & new_n5207;
  assign new_n11802 = ~new_n11800 & ~new_n11801;
  assign new_n11803 = ~new_n5243 & ~new_n11802;
  assign new_n11804 = ~new_n5207 & n3788;
  assign new_n11805 = n3820 & new_n5207;
  assign new_n11806 = ~new_n11804 & ~new_n11805;
  assign new_n11807 = ~new_n11806 & new_n5243;
  assign new_n11808 = ~new_n11803 & ~new_n11807;
  assign new_n11809 = ~new_n11808 & new_n5170;
  assign new_n11810 = ~new_n11799 & ~new_n11809;
  assign new_n11811 = ~new_n5139 & ~new_n11810;
  assign new_n11812 = ~new_n5207 & n3852;
  assign new_n11813 = n3884 & new_n5207;
  assign new_n11814 = ~new_n11812 & ~new_n11813;
  assign new_n11815 = ~new_n5243 & ~new_n11814;
  assign new_n11816 = ~new_n5207 & n3916;
  assign new_n11817 = n3948 & new_n5207;
  assign new_n11818 = ~new_n11816 & ~new_n11817;
  assign new_n11819 = ~new_n11818 & new_n5243;
  assign new_n11820 = ~new_n11815 & ~new_n11819;
  assign new_n11821 = ~new_n5170 & ~new_n11820;
  assign new_n11822 = ~new_n5207 & n3980;
  assign new_n11823 = n4012 & new_n5207;
  assign new_n11824 = ~new_n11822 & ~new_n11823;
  assign new_n11825 = ~new_n5243 & ~new_n11824;
  assign new_n11826 = ~new_n5207 & n4044;
  assign new_n11827 = n4076 & new_n5207;
  assign new_n11828 = ~new_n11826 & ~new_n11827;
  assign new_n11829 = ~new_n11828 & new_n5243;
  assign new_n11830 = ~new_n11825 & ~new_n11829;
  assign new_n11831 = ~new_n11830 & new_n5170;
  assign new_n11832 = ~new_n11821 & ~new_n11831;
  assign new_n11833 = ~new_n11832 & new_n5139;
  assign new_n11834 = ~new_n11811 & ~new_n11833;
  assign new_n11835 = ~new_n11834 & new_n5011;
  assign new_n11836 = ~new_n11789 & ~new_n11835;
  assign new_n11837 = ~new_n11836 & new_n5031;
  assign new_n11838 = ~new_n11743 & ~new_n11837;
  assign new_n11839 = ~new_n5077 & ~new_n11838;
  assign new_n11840 = ~new_n5207 & n2076;
  assign new_n11841 = n2108 & new_n5207;
  assign new_n11842 = ~new_n11840 & ~new_n11841;
  assign new_n11843 = ~new_n5243 & ~new_n11842;
  assign new_n11844 = ~new_n5207 & n2140;
  assign new_n11845 = n2172 & new_n5207;
  assign new_n11846 = ~new_n11844 & ~new_n11845;
  assign new_n11847 = ~new_n11846 & new_n5243;
  assign new_n11848 = ~new_n11843 & ~new_n11847;
  assign new_n11849 = ~new_n5170 & ~new_n11848;
  assign new_n11850 = ~new_n5207 & n2204;
  assign new_n11851 = n2236 & new_n5207;
  assign new_n11852 = ~new_n11850 & ~new_n11851;
  assign new_n11853 = ~new_n5243 & ~new_n11852;
  assign new_n11854 = ~new_n5207 & n2268;
  assign new_n11855 = n2300 & new_n5207;
  assign new_n11856 = ~new_n11854 & ~new_n11855;
  assign new_n11857 = ~new_n11856 & new_n5243;
  assign new_n11858 = ~new_n11853 & ~new_n11857;
  assign new_n11859 = ~new_n11858 & new_n5170;
  assign new_n11860 = ~new_n11849 & ~new_n11859;
  assign new_n11861 = ~new_n5139 & ~new_n11860;
  assign new_n11862 = ~new_n5207 & n2332;
  assign new_n11863 = n2364 & new_n5207;
  assign new_n11864 = ~new_n11862 & ~new_n11863;
  assign new_n11865 = ~new_n5243 & ~new_n11864;
  assign new_n11866 = ~new_n5207 & n2396;
  assign new_n11867 = n2428 & new_n5207;
  assign new_n11868 = ~new_n11866 & ~new_n11867;
  assign new_n11869 = ~new_n11868 & new_n5243;
  assign new_n11870 = ~new_n11865 & ~new_n11869;
  assign new_n11871 = ~new_n5170 & ~new_n11870;
  assign new_n11872 = ~new_n5207 & n2460;
  assign new_n11873 = n2492 & new_n5207;
  assign new_n11874 = ~new_n11872 & ~new_n11873;
  assign new_n11875 = ~new_n5243 & ~new_n11874;
  assign new_n11876 = ~new_n5207 & n2524;
  assign new_n11877 = n2556 & new_n5207;
  assign new_n11878 = ~new_n11876 & ~new_n11877;
  assign new_n11879 = ~new_n11878 & new_n5243;
  assign new_n11880 = ~new_n11875 & ~new_n11879;
  assign new_n11881 = ~new_n11880 & new_n5170;
  assign new_n11882 = ~new_n11871 & ~new_n11881;
  assign new_n11883 = ~new_n11882 & new_n5139;
  assign new_n11884 = ~new_n11861 & ~new_n11883;
  assign new_n11885 = ~new_n5011 & ~new_n11884;
  assign new_n11886 = ~new_n5207 & n2588;
  assign new_n11887 = n2620 & new_n5207;
  assign new_n11888 = ~new_n11886 & ~new_n11887;
  assign new_n11889 = ~new_n5243 & ~new_n11888;
  assign new_n11890 = ~new_n5207 & n2652;
  assign new_n11891 = n2684 & new_n5207;
  assign new_n11892 = ~new_n11890 & ~new_n11891;
  assign new_n11893 = ~new_n11892 & new_n5243;
  assign new_n11894 = ~new_n11889 & ~new_n11893;
  assign new_n11895 = ~new_n5170 & ~new_n11894;
  assign new_n11896 = ~new_n5207 & n2716;
  assign new_n11897 = n2748 & new_n5207;
  assign new_n11898 = ~new_n11896 & ~new_n11897;
  assign new_n11899 = ~new_n5243 & ~new_n11898;
  assign new_n11900 = ~new_n5207 & n2780;
  assign new_n11901 = n2812 & new_n5207;
  assign new_n11902 = ~new_n11900 & ~new_n11901;
  assign new_n11903 = ~new_n11902 & new_n5243;
  assign new_n11904 = ~new_n11899 & ~new_n11903;
  assign new_n11905 = ~new_n11904 & new_n5170;
  assign new_n11906 = ~new_n11895 & ~new_n11905;
  assign new_n11907 = ~new_n5139 & ~new_n11906;
  assign new_n11908 = ~new_n5207 & n2844;
  assign new_n11909 = n2876 & new_n5207;
  assign new_n11910 = ~new_n11908 & ~new_n11909;
  assign new_n11911 = ~new_n5243 & ~new_n11910;
  assign new_n11912 = ~new_n5207 & n2908;
  assign new_n11913 = n2940 & new_n5207;
  assign new_n11914 = ~new_n11912 & ~new_n11913;
  assign new_n11915 = ~new_n11914 & new_n5243;
  assign new_n11916 = ~new_n11911 & ~new_n11915;
  assign new_n11917 = ~new_n5170 & ~new_n11916;
  assign new_n11918 = ~new_n5207 & n2972;
  assign new_n11919 = n3004 & new_n5207;
  assign new_n11920 = ~new_n11918 & ~new_n11919;
  assign new_n11921 = ~new_n5243 & ~new_n11920;
  assign new_n11922 = ~new_n5207 & n3036;
  assign new_n11923 = n3068 & new_n5207;
  assign new_n11924 = ~new_n11922 & ~new_n11923;
  assign new_n11925 = ~new_n11924 & new_n5243;
  assign new_n11926 = ~new_n11921 & ~new_n11925;
  assign new_n11927 = ~new_n11926 & new_n5170;
  assign new_n11928 = ~new_n11917 & ~new_n11927;
  assign new_n11929 = ~new_n11928 & new_n5139;
  assign new_n11930 = ~new_n11907 & ~new_n11929;
  assign new_n11931 = ~new_n11930 & new_n5011;
  assign new_n11932 = ~new_n11885 & ~new_n11931;
  assign new_n11933 = ~new_n5031 & ~new_n11932;
  assign new_n11934 = ~new_n5207 & n3100;
  assign new_n11935 = n3132 & new_n5207;
  assign new_n11936 = ~new_n11934 & ~new_n11935;
  assign new_n11937 = ~new_n5243 & ~new_n11936;
  assign new_n11938 = ~new_n5207 & n3164;
  assign new_n11939 = n3196 & new_n5207;
  assign new_n11940 = ~new_n11938 & ~new_n11939;
  assign new_n11941 = ~new_n11940 & new_n5243;
  assign new_n11942 = ~new_n11937 & ~new_n11941;
  assign new_n11943 = ~new_n5170 & ~new_n11942;
  assign new_n11944 = ~new_n5207 & n3228;
  assign new_n11945 = n3260 & new_n5207;
  assign new_n11946 = ~new_n11944 & ~new_n11945;
  assign new_n11947 = ~new_n5243 & ~new_n11946;
  assign new_n11948 = ~new_n5207 & n3292;
  assign new_n11949 = n3324 & new_n5207;
  assign new_n11950 = ~new_n11948 & ~new_n11949;
  assign new_n11951 = ~new_n11950 & new_n5243;
  assign new_n11952 = ~new_n11947 & ~new_n11951;
  assign new_n11953 = ~new_n11952 & new_n5170;
  assign new_n11954 = ~new_n11943 & ~new_n11953;
  assign new_n11955 = ~new_n5139 & ~new_n11954;
  assign new_n11956 = ~new_n5207 & n3356;
  assign new_n11957 = n3388 & new_n5207;
  assign new_n11958 = ~new_n11956 & ~new_n11957;
  assign new_n11959 = ~new_n5243 & ~new_n11958;
  assign new_n11960 = ~new_n5207 & n3420;
  assign new_n11961 = n3452 & new_n5207;
  assign new_n11962 = ~new_n11960 & ~new_n11961;
  assign new_n11963 = ~new_n11962 & new_n5243;
  assign new_n11964 = ~new_n11959 & ~new_n11963;
  assign new_n11965 = ~new_n5170 & ~new_n11964;
  assign new_n11966 = ~new_n5207 & n3484;
  assign new_n11967 = n3516 & new_n5207;
  assign new_n11968 = ~new_n11966 & ~new_n11967;
  assign new_n11969 = ~new_n5243 & ~new_n11968;
  assign new_n11970 = ~new_n5207 & n3548;
  assign new_n11971 = n3580 & new_n5207;
  assign new_n11972 = ~new_n11970 & ~new_n11971;
  assign new_n11973 = ~new_n11972 & new_n5243;
  assign new_n11974 = ~new_n11969 & ~new_n11973;
  assign new_n11975 = ~new_n11974 & new_n5170;
  assign new_n11976 = ~new_n11965 & ~new_n11975;
  assign new_n11977 = ~new_n11976 & new_n5139;
  assign new_n11978 = ~new_n11955 & ~new_n11977;
  assign new_n11979 = ~new_n5011 & ~new_n11978;
  assign new_n11980 = ~new_n5207 & n3612;
  assign new_n11981 = n3644 & new_n5207;
  assign new_n11982 = ~new_n11980 & ~new_n11981;
  assign new_n11983 = ~new_n5243 & ~new_n11982;
  assign new_n11984 = ~new_n5207 & n3676;
  assign new_n11985 = n3708 & new_n5207;
  assign new_n11986 = ~new_n11984 & ~new_n11985;
  assign new_n11987 = ~new_n11986 & new_n5243;
  assign new_n11988 = ~new_n11983 & ~new_n11987;
  assign new_n11989 = ~new_n5170 & ~new_n11988;
  assign new_n11990 = ~new_n5207 & n3740;
  assign new_n11991 = n3772 & new_n5207;
  assign new_n11992 = ~new_n11990 & ~new_n11991;
  assign new_n11993 = ~new_n5243 & ~new_n11992;
  assign new_n11994 = ~new_n5207 & n3804;
  assign new_n11995 = n3836 & new_n5207;
  assign new_n11996 = ~new_n11994 & ~new_n11995;
  assign new_n11997 = ~new_n11996 & new_n5243;
  assign new_n11998 = ~new_n11993 & ~new_n11997;
  assign new_n11999 = ~new_n11998 & new_n5170;
  assign new_n12000 = ~new_n11989 & ~new_n11999;
  assign new_n12001 = ~new_n5139 & ~new_n12000;
  assign new_n12002 = ~new_n5207 & n3868;
  assign new_n12003 = n3900 & new_n5207;
  assign new_n12004 = ~new_n12002 & ~new_n12003;
  assign new_n12005 = ~new_n5243 & ~new_n12004;
  assign new_n12006 = ~new_n5207 & n3932;
  assign new_n12007 = n3964 & new_n5207;
  assign new_n12008 = ~new_n12006 & ~new_n12007;
  assign new_n12009 = ~new_n12008 & new_n5243;
  assign new_n12010 = ~new_n12005 & ~new_n12009;
  assign new_n12011 = ~new_n5170 & ~new_n12010;
  assign new_n12012 = ~new_n5207 & n3996;
  assign new_n12013 = n4028 & new_n5207;
  assign new_n12014 = ~new_n12012 & ~new_n12013;
  assign new_n12015 = ~new_n5243 & ~new_n12014;
  assign new_n12016 = ~new_n5207 & n4060;
  assign new_n12017 = n4092 & new_n5207;
  assign new_n12018 = ~new_n12016 & ~new_n12017;
  assign new_n12019 = ~new_n12018 & new_n5243;
  assign new_n12020 = ~new_n12015 & ~new_n12019;
  assign new_n12021 = ~new_n12020 & new_n5170;
  assign new_n12022 = ~new_n12011 & ~new_n12021;
  assign new_n12023 = ~new_n12022 & new_n5139;
  assign new_n12024 = ~new_n12001 & ~new_n12023;
  assign new_n12025 = ~new_n12024 & new_n5011;
  assign new_n12026 = ~new_n11979 & ~new_n12025;
  assign new_n12027 = ~new_n12026 & new_n5031;
  assign new_n12028 = ~new_n11933 & ~new_n12027;
  assign new_n12029 = ~new_n12028 & new_n5077;
  assign new_n12030 = ~new_n11839 & ~new_n12029;
  assign new_n12031 = ~new_n12030 & new_n8902;
  assign new_n12032 = ~new_n5207 & n2052;
  assign new_n12033 = n2084 & new_n5207;
  assign new_n12034 = ~new_n12032 & ~new_n12033;
  assign new_n12035 = ~new_n5243 & ~new_n12034;
  assign new_n12036 = ~new_n5207 & n2116;
  assign new_n12037 = n2148 & new_n5207;
  assign new_n12038 = ~new_n12036 & ~new_n12037;
  assign new_n12039 = ~new_n12038 & new_n5243;
  assign new_n12040 = ~new_n12035 & ~new_n12039;
  assign new_n12041 = ~new_n5170 & ~new_n12040;
  assign new_n12042 = ~new_n5207 & n2180;
  assign new_n12043 = n2212 & new_n5207;
  assign new_n12044 = ~new_n12042 & ~new_n12043;
  assign new_n12045 = ~new_n5243 & ~new_n12044;
  assign new_n12046 = ~new_n5207 & n2244;
  assign new_n12047 = n2276 & new_n5207;
  assign new_n12048 = ~new_n12046 & ~new_n12047;
  assign new_n12049 = ~new_n12048 & new_n5243;
  assign new_n12050 = ~new_n12045 & ~new_n12049;
  assign new_n12051 = ~new_n12050 & new_n5170;
  assign new_n12052 = ~new_n12041 & ~new_n12051;
  assign new_n12053 = ~new_n5139 & ~new_n12052;
  assign new_n12054 = ~new_n5207 & n2308;
  assign new_n12055 = n2340 & new_n5207;
  assign new_n12056 = ~new_n12054 & ~new_n12055;
  assign new_n12057 = ~new_n5243 & ~new_n12056;
  assign new_n12058 = ~new_n5207 & n2372;
  assign new_n12059 = n2404 & new_n5207;
  assign new_n12060 = ~new_n12058 & ~new_n12059;
  assign new_n12061 = ~new_n12060 & new_n5243;
  assign new_n12062 = ~new_n12057 & ~new_n12061;
  assign new_n12063 = ~new_n5170 & ~new_n12062;
  assign new_n12064 = ~new_n5207 & n2436;
  assign new_n12065 = n2468 & new_n5207;
  assign new_n12066 = ~new_n12064 & ~new_n12065;
  assign new_n12067 = ~new_n5243 & ~new_n12066;
  assign new_n12068 = ~new_n5207 & n2500;
  assign new_n12069 = n2532 & new_n5207;
  assign new_n12070 = ~new_n12068 & ~new_n12069;
  assign new_n12071 = ~new_n12070 & new_n5243;
  assign new_n12072 = ~new_n12067 & ~new_n12071;
  assign new_n12073 = ~new_n12072 & new_n5170;
  assign new_n12074 = ~new_n12063 & ~new_n12073;
  assign new_n12075 = ~new_n12074 & new_n5139;
  assign new_n12076 = ~new_n12053 & ~new_n12075;
  assign new_n12077 = ~new_n5011 & ~new_n12076;
  assign new_n12078 = ~new_n5207 & n2564;
  assign new_n12079 = n2596 & new_n5207;
  assign new_n12080 = ~new_n12078 & ~new_n12079;
  assign new_n12081 = ~new_n5243 & ~new_n12080;
  assign new_n12082 = ~new_n5207 & n2628;
  assign new_n12083 = n2660 & new_n5207;
  assign new_n12084 = ~new_n12082 & ~new_n12083;
  assign new_n12085 = ~new_n12084 & new_n5243;
  assign new_n12086 = ~new_n12081 & ~new_n12085;
  assign new_n12087 = ~new_n5170 & ~new_n12086;
  assign new_n12088 = ~new_n5207 & n2692;
  assign new_n12089 = n2724 & new_n5207;
  assign new_n12090 = ~new_n12088 & ~new_n12089;
  assign new_n12091 = ~new_n5243 & ~new_n12090;
  assign new_n12092 = ~new_n5207 & n2756;
  assign new_n12093 = n2788 & new_n5207;
  assign new_n12094 = ~new_n12092 & ~new_n12093;
  assign new_n12095 = ~new_n12094 & new_n5243;
  assign new_n12096 = ~new_n12091 & ~new_n12095;
  assign new_n12097 = ~new_n12096 & new_n5170;
  assign new_n12098 = ~new_n12087 & ~new_n12097;
  assign new_n12099 = ~new_n5139 & ~new_n12098;
  assign new_n12100 = ~new_n5207 & n2820;
  assign new_n12101 = n2852 & new_n5207;
  assign new_n12102 = ~new_n12100 & ~new_n12101;
  assign new_n12103 = ~new_n5243 & ~new_n12102;
  assign new_n12104 = ~new_n5207 & n2884;
  assign new_n12105 = n2916 & new_n5207;
  assign new_n12106 = ~new_n12104 & ~new_n12105;
  assign new_n12107 = ~new_n12106 & new_n5243;
  assign new_n12108 = ~new_n12103 & ~new_n12107;
  assign new_n12109 = ~new_n5170 & ~new_n12108;
  assign new_n12110 = ~new_n5207 & n2948;
  assign new_n12111 = n2980 & new_n5207;
  assign new_n12112 = ~new_n12110 & ~new_n12111;
  assign new_n12113 = ~new_n5243 & ~new_n12112;
  assign new_n12114 = ~new_n5207 & n3012;
  assign new_n12115 = n3044 & new_n5207;
  assign new_n12116 = ~new_n12114 & ~new_n12115;
  assign new_n12117 = ~new_n12116 & new_n5243;
  assign new_n12118 = ~new_n12113 & ~new_n12117;
  assign new_n12119 = ~new_n12118 & new_n5170;
  assign new_n12120 = ~new_n12109 & ~new_n12119;
  assign new_n12121 = ~new_n12120 & new_n5139;
  assign new_n12122 = ~new_n12099 & ~new_n12121;
  assign new_n12123 = ~new_n12122 & new_n5011;
  assign new_n12124 = ~new_n12077 & ~new_n12123;
  assign new_n12125 = ~new_n5031 & ~new_n12124;
  assign new_n12126 = ~new_n5207 & n3076;
  assign new_n12127 = n3108 & new_n5207;
  assign new_n12128 = ~new_n12126 & ~new_n12127;
  assign new_n12129 = ~new_n5243 & ~new_n12128;
  assign new_n12130 = ~new_n5207 & n3140;
  assign new_n12131 = n3172 & new_n5207;
  assign new_n12132 = ~new_n12130 & ~new_n12131;
  assign new_n12133 = ~new_n12132 & new_n5243;
  assign new_n12134 = ~new_n12129 & ~new_n12133;
  assign new_n12135 = ~new_n5170 & ~new_n12134;
  assign new_n12136 = ~new_n5207 & n3204;
  assign new_n12137 = n3236 & new_n5207;
  assign new_n12138 = ~new_n12136 & ~new_n12137;
  assign new_n12139 = ~new_n5243 & ~new_n12138;
  assign new_n12140 = ~new_n5207 & n3268;
  assign new_n12141 = n3300 & new_n5207;
  assign new_n12142 = ~new_n12140 & ~new_n12141;
  assign new_n12143 = ~new_n12142 & new_n5243;
  assign new_n12144 = ~new_n12139 & ~new_n12143;
  assign new_n12145 = ~new_n12144 & new_n5170;
  assign new_n12146 = ~new_n12135 & ~new_n12145;
  assign new_n12147 = ~new_n5139 & ~new_n12146;
  assign new_n12148 = ~new_n5207 & n3332;
  assign new_n12149 = n3364 & new_n5207;
  assign new_n12150 = ~new_n12148 & ~new_n12149;
  assign new_n12151 = ~new_n5243 & ~new_n12150;
  assign new_n12152 = ~new_n5207 & n3396;
  assign new_n12153 = n3428 & new_n5207;
  assign new_n12154 = ~new_n12152 & ~new_n12153;
  assign new_n12155 = ~new_n12154 & new_n5243;
  assign new_n12156 = ~new_n12151 & ~new_n12155;
  assign new_n12157 = ~new_n5170 & ~new_n12156;
  assign new_n12158 = ~new_n5207 & n3460;
  assign new_n12159 = n3492 & new_n5207;
  assign new_n12160 = ~new_n12158 & ~new_n12159;
  assign new_n12161 = ~new_n5243 & ~new_n12160;
  assign new_n12162 = ~new_n5207 & n3524;
  assign new_n12163 = n3556 & new_n5207;
  assign new_n12164 = ~new_n12162 & ~new_n12163;
  assign new_n12165 = ~new_n12164 & new_n5243;
  assign new_n12166 = ~new_n12161 & ~new_n12165;
  assign new_n12167 = ~new_n12166 & new_n5170;
  assign new_n12168 = ~new_n12157 & ~new_n12167;
  assign new_n12169 = ~new_n12168 & new_n5139;
  assign new_n12170 = ~new_n12147 & ~new_n12169;
  assign new_n12171 = ~new_n5011 & ~new_n12170;
  assign new_n12172 = ~new_n5207 & n3588;
  assign new_n12173 = n3620 & new_n5207;
  assign new_n12174 = ~new_n12172 & ~new_n12173;
  assign new_n12175 = ~new_n5243 & ~new_n12174;
  assign new_n12176 = ~new_n5207 & n3652;
  assign new_n12177 = n3684 & new_n5207;
  assign new_n12178 = ~new_n12176 & ~new_n12177;
  assign new_n12179 = ~new_n12178 & new_n5243;
  assign new_n12180 = ~new_n12175 & ~new_n12179;
  assign new_n12181 = ~new_n5170 & ~new_n12180;
  assign new_n12182 = ~new_n5207 & n3716;
  assign new_n12183 = n3748 & new_n5207;
  assign new_n12184 = ~new_n12182 & ~new_n12183;
  assign new_n12185 = ~new_n5243 & ~new_n12184;
  assign new_n12186 = ~new_n5207 & n3780;
  assign new_n12187 = n3812 & new_n5207;
  assign new_n12188 = ~new_n12186 & ~new_n12187;
  assign new_n12189 = ~new_n12188 & new_n5243;
  assign new_n12190 = ~new_n12185 & ~new_n12189;
  assign new_n12191 = ~new_n12190 & new_n5170;
  assign new_n12192 = ~new_n12181 & ~new_n12191;
  assign new_n12193 = ~new_n5139 & ~new_n12192;
  assign new_n12194 = ~new_n5207 & n3844;
  assign new_n12195 = n3876 & new_n5207;
  assign new_n12196 = ~new_n12194 & ~new_n12195;
  assign new_n12197 = ~new_n5243 & ~new_n12196;
  assign new_n12198 = ~new_n5207 & n3908;
  assign new_n12199 = n3940 & new_n5207;
  assign new_n12200 = ~new_n12198 & ~new_n12199;
  assign new_n12201 = ~new_n12200 & new_n5243;
  assign new_n12202 = ~new_n12197 & ~new_n12201;
  assign new_n12203 = ~new_n5170 & ~new_n12202;
  assign new_n12204 = ~new_n5207 & n3972;
  assign new_n12205 = n4004 & new_n5207;
  assign new_n12206 = ~new_n12204 & ~new_n12205;
  assign new_n12207 = ~new_n5243 & ~new_n12206;
  assign new_n12208 = ~new_n5207 & n4036;
  assign new_n12209 = n4068 & new_n5207;
  assign new_n12210 = ~new_n12208 & ~new_n12209;
  assign new_n12211 = ~new_n12210 & new_n5243;
  assign new_n12212 = ~new_n12207 & ~new_n12211;
  assign new_n12213 = ~new_n12212 & new_n5170;
  assign new_n12214 = ~new_n12203 & ~new_n12213;
  assign new_n12215 = ~new_n12214 & new_n5139;
  assign new_n12216 = ~new_n12193 & ~new_n12215;
  assign new_n12217 = ~new_n12216 & new_n5011;
  assign new_n12218 = ~new_n12171 & ~new_n12217;
  assign new_n12219 = ~new_n12218 & new_n5031;
  assign new_n12220 = ~new_n12125 & ~new_n12219;
  assign new_n12221 = ~new_n12220 & new_n5114;
  assign new_n12222 = ~new_n5462 & ~new_n11838;
  assign new_n12223 = ~new_n12221 & ~new_n12222;
  assign new_n12224 = ~new_n5207 & n2068;
  assign new_n12225 = n2100 & new_n5207;
  assign new_n12226 = ~new_n12224 & ~new_n12225;
  assign new_n12227 = ~new_n5243 & ~new_n12226;
  assign new_n12228 = ~new_n5207 & n2132;
  assign new_n12229 = n2164 & new_n5207;
  assign new_n12230 = ~new_n12228 & ~new_n12229;
  assign new_n12231 = ~new_n12230 & new_n5243;
  assign new_n12232 = ~new_n12227 & ~new_n12231;
  assign new_n12233 = ~new_n5170 & ~new_n12232;
  assign new_n12234 = ~new_n5207 & n2196;
  assign new_n12235 = n2228 & new_n5207;
  assign new_n12236 = ~new_n12234 & ~new_n12235;
  assign new_n12237 = ~new_n5243 & ~new_n12236;
  assign new_n12238 = ~new_n5207 & n2260;
  assign new_n12239 = n2292 & new_n5207;
  assign new_n12240 = ~new_n12238 & ~new_n12239;
  assign new_n12241 = ~new_n12240 & new_n5243;
  assign new_n12242 = ~new_n12237 & ~new_n12241;
  assign new_n12243 = ~new_n12242 & new_n5170;
  assign new_n12244 = ~new_n12233 & ~new_n12243;
  assign new_n12245 = ~new_n5139 & ~new_n12244;
  assign new_n12246 = ~new_n5207 & n2324;
  assign new_n12247 = n2356 & new_n5207;
  assign new_n12248 = ~new_n12246 & ~new_n12247;
  assign new_n12249 = ~new_n5243 & ~new_n12248;
  assign new_n12250 = ~new_n5207 & n2388;
  assign new_n12251 = n2420 & new_n5207;
  assign new_n12252 = ~new_n12250 & ~new_n12251;
  assign new_n12253 = ~new_n12252 & new_n5243;
  assign new_n12254 = ~new_n12249 & ~new_n12253;
  assign new_n12255 = ~new_n5170 & ~new_n12254;
  assign new_n12256 = ~new_n5207 & n2452;
  assign new_n12257 = n2484 & new_n5207;
  assign new_n12258 = ~new_n12256 & ~new_n12257;
  assign new_n12259 = ~new_n5243 & ~new_n12258;
  assign new_n12260 = ~new_n5207 & n2516;
  assign new_n12261 = n2548 & new_n5207;
  assign new_n12262 = ~new_n12260 & ~new_n12261;
  assign new_n12263 = ~new_n12262 & new_n5243;
  assign new_n12264 = ~new_n12259 & ~new_n12263;
  assign new_n12265 = ~new_n12264 & new_n5170;
  assign new_n12266 = ~new_n12255 & ~new_n12265;
  assign new_n12267 = ~new_n12266 & new_n5139;
  assign new_n12268 = ~new_n12245 & ~new_n12267;
  assign new_n12269 = ~new_n5011 & ~new_n12268;
  assign new_n12270 = ~new_n5207 & n2580;
  assign new_n12271 = n2612 & new_n5207;
  assign new_n12272 = ~new_n12270 & ~new_n12271;
  assign new_n12273 = ~new_n5243 & ~new_n12272;
  assign new_n12274 = ~new_n5207 & n2644;
  assign new_n12275 = n2676 & new_n5207;
  assign new_n12276 = ~new_n12274 & ~new_n12275;
  assign new_n12277 = ~new_n12276 & new_n5243;
  assign new_n12278 = ~new_n12273 & ~new_n12277;
  assign new_n12279 = ~new_n5170 & ~new_n12278;
  assign new_n12280 = ~new_n5207 & n2708;
  assign new_n12281 = n2740 & new_n5207;
  assign new_n12282 = ~new_n12280 & ~new_n12281;
  assign new_n12283 = ~new_n5243 & ~new_n12282;
  assign new_n12284 = ~new_n5207 & n2772;
  assign new_n12285 = n2804 & new_n5207;
  assign new_n12286 = ~new_n12284 & ~new_n12285;
  assign new_n12287 = ~new_n12286 & new_n5243;
  assign new_n12288 = ~new_n12283 & ~new_n12287;
  assign new_n12289 = ~new_n12288 & new_n5170;
  assign new_n12290 = ~new_n12279 & ~new_n12289;
  assign new_n12291 = ~new_n5139 & ~new_n12290;
  assign new_n12292 = ~new_n5207 & n2836;
  assign new_n12293 = n2868 & new_n5207;
  assign new_n12294 = ~new_n12292 & ~new_n12293;
  assign new_n12295 = ~new_n5243 & ~new_n12294;
  assign new_n12296 = ~new_n5207 & n2900;
  assign new_n12297 = n2932 & new_n5207;
  assign new_n12298 = ~new_n12296 & ~new_n12297;
  assign new_n12299 = ~new_n12298 & new_n5243;
  assign new_n12300 = ~new_n12295 & ~new_n12299;
  assign new_n12301 = ~new_n5170 & ~new_n12300;
  assign new_n12302 = ~new_n5207 & n2964;
  assign new_n12303 = n2996 & new_n5207;
  assign new_n12304 = ~new_n12302 & ~new_n12303;
  assign new_n12305 = ~new_n5243 & ~new_n12304;
  assign new_n12306 = ~new_n5207 & n3028;
  assign new_n12307 = n3060 & new_n5207;
  assign new_n12308 = ~new_n12306 & ~new_n12307;
  assign new_n12309 = ~new_n12308 & new_n5243;
  assign new_n12310 = ~new_n12305 & ~new_n12309;
  assign new_n12311 = ~new_n12310 & new_n5170;
  assign new_n12312 = ~new_n12301 & ~new_n12311;
  assign new_n12313 = ~new_n12312 & new_n5139;
  assign new_n12314 = ~new_n12291 & ~new_n12313;
  assign new_n12315 = ~new_n12314 & new_n5011;
  assign new_n12316 = ~new_n12269 & ~new_n12315;
  assign new_n12317 = ~new_n5031 & ~new_n12316;
  assign new_n12318 = ~new_n5207 & n3092;
  assign new_n12319 = n3124 & new_n5207;
  assign new_n12320 = ~new_n12318 & ~new_n12319;
  assign new_n12321 = ~new_n5243 & ~new_n12320;
  assign new_n12322 = ~new_n5207 & n3156;
  assign new_n12323 = n3188 & new_n5207;
  assign new_n12324 = ~new_n12322 & ~new_n12323;
  assign new_n12325 = ~new_n12324 & new_n5243;
  assign new_n12326 = ~new_n12321 & ~new_n12325;
  assign new_n12327 = ~new_n5170 & ~new_n12326;
  assign new_n12328 = ~new_n5207 & n3220;
  assign new_n12329 = n3252 & new_n5207;
  assign new_n12330 = ~new_n12328 & ~new_n12329;
  assign new_n12331 = ~new_n5243 & ~new_n12330;
  assign new_n12332 = ~new_n5207 & n3284;
  assign new_n12333 = n3316 & new_n5207;
  assign new_n12334 = ~new_n12332 & ~new_n12333;
  assign new_n12335 = ~new_n12334 & new_n5243;
  assign new_n12336 = ~new_n12331 & ~new_n12335;
  assign new_n12337 = ~new_n12336 & new_n5170;
  assign new_n12338 = ~new_n12327 & ~new_n12337;
  assign new_n12339 = ~new_n5139 & ~new_n12338;
  assign new_n12340 = ~new_n5207 & n3348;
  assign new_n12341 = n3380 & new_n5207;
  assign new_n12342 = ~new_n12340 & ~new_n12341;
  assign new_n12343 = ~new_n5243 & ~new_n12342;
  assign new_n12344 = ~new_n5207 & n3412;
  assign new_n12345 = n3444 & new_n5207;
  assign new_n12346 = ~new_n12344 & ~new_n12345;
  assign new_n12347 = ~new_n12346 & new_n5243;
  assign new_n12348 = ~new_n12343 & ~new_n12347;
  assign new_n12349 = ~new_n5170 & ~new_n12348;
  assign new_n12350 = ~new_n5207 & n3476;
  assign new_n12351 = n3508 & new_n5207;
  assign new_n12352 = ~new_n12350 & ~new_n12351;
  assign new_n12353 = ~new_n5243 & ~new_n12352;
  assign new_n12354 = ~new_n5207 & n3540;
  assign new_n12355 = n3572 & new_n5207;
  assign new_n12356 = ~new_n12354 & ~new_n12355;
  assign new_n12357 = ~new_n12356 & new_n5243;
  assign new_n12358 = ~new_n12353 & ~new_n12357;
  assign new_n12359 = ~new_n12358 & new_n5170;
  assign new_n12360 = ~new_n12349 & ~new_n12359;
  assign new_n12361 = ~new_n12360 & new_n5139;
  assign new_n12362 = ~new_n12339 & ~new_n12361;
  assign new_n12363 = ~new_n5011 & ~new_n12362;
  assign new_n12364 = ~new_n5207 & n3604;
  assign new_n12365 = n3636 & new_n5207;
  assign new_n12366 = ~new_n12364 & ~new_n12365;
  assign new_n12367 = ~new_n5243 & ~new_n12366;
  assign new_n12368 = ~new_n5207 & n3668;
  assign new_n12369 = n3700 & new_n5207;
  assign new_n12370 = ~new_n12368 & ~new_n12369;
  assign new_n12371 = ~new_n12370 & new_n5243;
  assign new_n12372 = ~new_n12367 & ~new_n12371;
  assign new_n12373 = ~new_n5170 & ~new_n12372;
  assign new_n12374 = ~new_n5207 & n3732;
  assign new_n12375 = n3764 & new_n5207;
  assign new_n12376 = ~new_n12374 & ~new_n12375;
  assign new_n12377 = ~new_n5243 & ~new_n12376;
  assign new_n12378 = ~new_n5207 & n3796;
  assign new_n12379 = n3828 & new_n5207;
  assign new_n12380 = ~new_n12378 & ~new_n12379;
  assign new_n12381 = ~new_n12380 & new_n5243;
  assign new_n12382 = ~new_n12377 & ~new_n12381;
  assign new_n12383 = ~new_n12382 & new_n5170;
  assign new_n12384 = ~new_n12373 & ~new_n12383;
  assign new_n12385 = ~new_n5139 & ~new_n12384;
  assign new_n12386 = ~new_n5207 & n3860;
  assign new_n12387 = n3892 & new_n5207;
  assign new_n12388 = ~new_n12386 & ~new_n12387;
  assign new_n12389 = ~new_n5243 & ~new_n12388;
  assign new_n12390 = ~new_n5207 & n3924;
  assign new_n12391 = n3956 & new_n5207;
  assign new_n12392 = ~new_n12390 & ~new_n12391;
  assign new_n12393 = ~new_n12392 & new_n5243;
  assign new_n12394 = ~new_n12389 & ~new_n12393;
  assign new_n12395 = ~new_n5170 & ~new_n12394;
  assign new_n12396 = ~new_n5207 & n3988;
  assign new_n12397 = n4020 & new_n5207;
  assign new_n12398 = ~new_n12396 & ~new_n12397;
  assign new_n12399 = ~new_n5243 & ~new_n12398;
  assign new_n12400 = ~new_n5207 & n4052;
  assign new_n12401 = n4084 & new_n5207;
  assign new_n12402 = ~new_n12400 & ~new_n12401;
  assign new_n12403 = ~new_n12402 & new_n5243;
  assign new_n12404 = ~new_n12399 & ~new_n12403;
  assign new_n12405 = ~new_n12404 & new_n5170;
  assign new_n12406 = ~new_n12395 & ~new_n12405;
  assign new_n12407 = ~new_n12406 & new_n5139;
  assign new_n12408 = ~new_n12385 & ~new_n12407;
  assign new_n12409 = ~new_n12408 & new_n5011;
  assign new_n12410 = ~new_n12363 & ~new_n12409;
  assign new_n12411 = ~new_n12410 & new_n5031;
  assign new_n12412 = ~new_n12317 & ~new_n12411;
  assign new_n12413 = ~new_n5115 & ~new_n12412;
  assign new_n12414 = ~new_n5116 & ~new_n12028;
  assign new_n12415 = ~new_n12413 & ~new_n12414;
  assign new_n12416 = new_n12223 & new_n12415;
  assign new_n12417 = ~new_n9289 & ~new_n12416;
  assign new_n12418 = ~new_n12031 & ~new_n12417;
  assign new_n12419 = ~new_n12416 & new_n8900;
  assign new_n12420 = ~new_n12030 & new_n8901;
  assign new_n12421 = ~new_n12419 & ~new_n12420;
  assign new_n12422 = ~new_n12028 & new_n4150;
  assign new_n12423 = ~new_n5170 & ~new_n9302;
  assign new_n12424 = ~new_n12422 & ~new_n12423;
  assign new_n12425 = new_n12421 & new_n12424;
  assign new_n12426 = new_n12418 & new_n12425;
  assign new_n12427 = ~new_n12426 & new_n8515;
  assign new_n12428 = ~new_n5207 & n2059;
  assign new_n12429 = n2091 & new_n5207;
  assign new_n12430 = ~new_n12428 & ~new_n12429;
  assign new_n12431 = ~new_n5243 & ~new_n12430;
  assign new_n12432 = ~new_n5207 & n2123;
  assign new_n12433 = n2155 & new_n5207;
  assign new_n12434 = ~new_n12432 & ~new_n12433;
  assign new_n12435 = ~new_n12434 & new_n5243;
  assign new_n12436 = ~new_n12431 & ~new_n12435;
  assign new_n12437 = ~new_n5170 & ~new_n12436;
  assign new_n12438 = ~new_n5207 & n2187;
  assign new_n12439 = n2219 & new_n5207;
  assign new_n12440 = ~new_n12438 & ~new_n12439;
  assign new_n12441 = ~new_n5243 & ~new_n12440;
  assign new_n12442 = ~new_n5207 & n2251;
  assign new_n12443 = n2283 & new_n5207;
  assign new_n12444 = ~new_n12442 & ~new_n12443;
  assign new_n12445 = ~new_n12444 & new_n5243;
  assign new_n12446 = ~new_n12441 & ~new_n12445;
  assign new_n12447 = ~new_n12446 & new_n5170;
  assign new_n12448 = ~new_n12437 & ~new_n12447;
  assign new_n12449 = ~new_n5139 & ~new_n12448;
  assign new_n12450 = ~new_n5207 & n2315;
  assign new_n12451 = n2347 & new_n5207;
  assign new_n12452 = ~new_n12450 & ~new_n12451;
  assign new_n12453 = ~new_n5243 & ~new_n12452;
  assign new_n12454 = ~new_n5207 & n2379;
  assign new_n12455 = n2411 & new_n5207;
  assign new_n12456 = ~new_n12454 & ~new_n12455;
  assign new_n12457 = ~new_n12456 & new_n5243;
  assign new_n12458 = ~new_n12453 & ~new_n12457;
  assign new_n12459 = ~new_n5170 & ~new_n12458;
  assign new_n12460 = ~new_n5207 & n2443;
  assign new_n12461 = n2475 & new_n5207;
  assign new_n12462 = ~new_n12460 & ~new_n12461;
  assign new_n12463 = ~new_n5243 & ~new_n12462;
  assign new_n12464 = ~new_n5207 & n2507;
  assign new_n12465 = n2539 & new_n5207;
  assign new_n12466 = ~new_n12464 & ~new_n12465;
  assign new_n12467 = ~new_n12466 & new_n5243;
  assign new_n12468 = ~new_n12463 & ~new_n12467;
  assign new_n12469 = ~new_n12468 & new_n5170;
  assign new_n12470 = ~new_n12459 & ~new_n12469;
  assign new_n12471 = ~new_n12470 & new_n5139;
  assign new_n12472 = ~new_n12449 & ~new_n12471;
  assign new_n12473 = ~new_n5011 & ~new_n12472;
  assign new_n12474 = ~new_n5207 & n2571;
  assign new_n12475 = n2603 & new_n5207;
  assign new_n12476 = ~new_n12474 & ~new_n12475;
  assign new_n12477 = ~new_n5243 & ~new_n12476;
  assign new_n12478 = ~new_n5207 & n2635;
  assign new_n12479 = n2667 & new_n5207;
  assign new_n12480 = ~new_n12478 & ~new_n12479;
  assign new_n12481 = ~new_n12480 & new_n5243;
  assign new_n12482 = ~new_n12477 & ~new_n12481;
  assign new_n12483 = ~new_n5170 & ~new_n12482;
  assign new_n12484 = ~new_n5207 & n2699;
  assign new_n12485 = n2731 & new_n5207;
  assign new_n12486 = ~new_n12484 & ~new_n12485;
  assign new_n12487 = ~new_n5243 & ~new_n12486;
  assign new_n12488 = ~new_n5207 & n2763;
  assign new_n12489 = n2795 & new_n5207;
  assign new_n12490 = ~new_n12488 & ~new_n12489;
  assign new_n12491 = ~new_n12490 & new_n5243;
  assign new_n12492 = ~new_n12487 & ~new_n12491;
  assign new_n12493 = ~new_n12492 & new_n5170;
  assign new_n12494 = ~new_n12483 & ~new_n12493;
  assign new_n12495 = ~new_n5139 & ~new_n12494;
  assign new_n12496 = ~new_n5207 & n2827;
  assign new_n12497 = n2859 & new_n5207;
  assign new_n12498 = ~new_n12496 & ~new_n12497;
  assign new_n12499 = ~new_n5243 & ~new_n12498;
  assign new_n12500 = ~new_n5207 & n2891;
  assign new_n12501 = n2923 & new_n5207;
  assign new_n12502 = ~new_n12500 & ~new_n12501;
  assign new_n12503 = ~new_n12502 & new_n5243;
  assign new_n12504 = ~new_n12499 & ~new_n12503;
  assign new_n12505 = ~new_n5170 & ~new_n12504;
  assign new_n12506 = ~new_n5207 & n2955;
  assign new_n12507 = n2987 & new_n5207;
  assign new_n12508 = ~new_n12506 & ~new_n12507;
  assign new_n12509 = ~new_n5243 & ~new_n12508;
  assign new_n12510 = ~new_n5207 & n3019;
  assign new_n12511 = n3051 & new_n5207;
  assign new_n12512 = ~new_n12510 & ~new_n12511;
  assign new_n12513 = ~new_n12512 & new_n5243;
  assign new_n12514 = ~new_n12509 & ~new_n12513;
  assign new_n12515 = ~new_n12514 & new_n5170;
  assign new_n12516 = ~new_n12505 & ~new_n12515;
  assign new_n12517 = ~new_n12516 & new_n5139;
  assign new_n12518 = ~new_n12495 & ~new_n12517;
  assign new_n12519 = ~new_n12518 & new_n5011;
  assign new_n12520 = ~new_n12473 & ~new_n12519;
  assign new_n12521 = ~new_n5031 & ~new_n12520;
  assign new_n12522 = ~new_n5207 & n3083;
  assign new_n12523 = n3115 & new_n5207;
  assign new_n12524 = ~new_n12522 & ~new_n12523;
  assign new_n12525 = ~new_n5243 & ~new_n12524;
  assign new_n12526 = ~new_n5207 & n3147;
  assign new_n12527 = n3179 & new_n5207;
  assign new_n12528 = ~new_n12526 & ~new_n12527;
  assign new_n12529 = ~new_n12528 & new_n5243;
  assign new_n12530 = ~new_n12525 & ~new_n12529;
  assign new_n12531 = ~new_n5170 & ~new_n12530;
  assign new_n12532 = ~new_n5207 & n3211;
  assign new_n12533 = n3243 & new_n5207;
  assign new_n12534 = ~new_n12532 & ~new_n12533;
  assign new_n12535 = ~new_n5243 & ~new_n12534;
  assign new_n12536 = ~new_n5207 & n3275;
  assign new_n12537 = n3307 & new_n5207;
  assign new_n12538 = ~new_n12536 & ~new_n12537;
  assign new_n12539 = ~new_n12538 & new_n5243;
  assign new_n12540 = ~new_n12535 & ~new_n12539;
  assign new_n12541 = ~new_n12540 & new_n5170;
  assign new_n12542 = ~new_n12531 & ~new_n12541;
  assign new_n12543 = ~new_n5139 & ~new_n12542;
  assign new_n12544 = ~new_n5207 & n3339;
  assign new_n12545 = n3371 & new_n5207;
  assign new_n12546 = ~new_n12544 & ~new_n12545;
  assign new_n12547 = ~new_n5243 & ~new_n12546;
  assign new_n12548 = ~new_n5207 & n3403;
  assign new_n12549 = n3435 & new_n5207;
  assign new_n12550 = ~new_n12548 & ~new_n12549;
  assign new_n12551 = ~new_n12550 & new_n5243;
  assign new_n12552 = ~new_n12547 & ~new_n12551;
  assign new_n12553 = ~new_n5170 & ~new_n12552;
  assign new_n12554 = ~new_n5207 & n3467;
  assign new_n12555 = n3499 & new_n5207;
  assign new_n12556 = ~new_n12554 & ~new_n12555;
  assign new_n12557 = ~new_n5243 & ~new_n12556;
  assign new_n12558 = ~new_n5207 & n3531;
  assign new_n12559 = n3563 & new_n5207;
  assign new_n12560 = ~new_n12558 & ~new_n12559;
  assign new_n12561 = ~new_n12560 & new_n5243;
  assign new_n12562 = ~new_n12557 & ~new_n12561;
  assign new_n12563 = ~new_n12562 & new_n5170;
  assign new_n12564 = ~new_n12553 & ~new_n12563;
  assign new_n12565 = ~new_n12564 & new_n5139;
  assign new_n12566 = ~new_n12543 & ~new_n12565;
  assign new_n12567 = ~new_n5011 & ~new_n12566;
  assign new_n12568 = ~new_n5207 & n3595;
  assign new_n12569 = n3627 & new_n5207;
  assign new_n12570 = ~new_n12568 & ~new_n12569;
  assign new_n12571 = ~new_n5243 & ~new_n12570;
  assign new_n12572 = ~new_n5207 & n3659;
  assign new_n12573 = n3691 & new_n5207;
  assign new_n12574 = ~new_n12572 & ~new_n12573;
  assign new_n12575 = ~new_n12574 & new_n5243;
  assign new_n12576 = ~new_n12571 & ~new_n12575;
  assign new_n12577 = ~new_n5170 & ~new_n12576;
  assign new_n12578 = ~new_n5207 & n3723;
  assign new_n12579 = n3755 & new_n5207;
  assign new_n12580 = ~new_n12578 & ~new_n12579;
  assign new_n12581 = ~new_n5243 & ~new_n12580;
  assign new_n12582 = ~new_n5207 & n3787;
  assign new_n12583 = n3819 & new_n5207;
  assign new_n12584 = ~new_n12582 & ~new_n12583;
  assign new_n12585 = ~new_n12584 & new_n5243;
  assign new_n12586 = ~new_n12581 & ~new_n12585;
  assign new_n12587 = ~new_n12586 & new_n5170;
  assign new_n12588 = ~new_n12577 & ~new_n12587;
  assign new_n12589 = ~new_n5139 & ~new_n12588;
  assign new_n12590 = ~new_n5207 & n3851;
  assign new_n12591 = n3883 & new_n5207;
  assign new_n12592 = ~new_n12590 & ~new_n12591;
  assign new_n12593 = ~new_n5243 & ~new_n12592;
  assign new_n12594 = ~new_n5207 & n3915;
  assign new_n12595 = n3947 & new_n5207;
  assign new_n12596 = ~new_n12594 & ~new_n12595;
  assign new_n12597 = ~new_n12596 & new_n5243;
  assign new_n12598 = ~new_n12593 & ~new_n12597;
  assign new_n12599 = ~new_n5170 & ~new_n12598;
  assign new_n12600 = ~new_n5207 & n3979;
  assign new_n12601 = n4011 & new_n5207;
  assign new_n12602 = ~new_n12600 & ~new_n12601;
  assign new_n12603 = ~new_n5243 & ~new_n12602;
  assign new_n12604 = ~new_n5207 & n4043;
  assign new_n12605 = n4075 & new_n5207;
  assign new_n12606 = ~new_n12604 & ~new_n12605;
  assign new_n12607 = ~new_n12606 & new_n5243;
  assign new_n12608 = ~new_n12603 & ~new_n12607;
  assign new_n12609 = ~new_n12608 & new_n5170;
  assign new_n12610 = ~new_n12599 & ~new_n12609;
  assign new_n12611 = ~new_n12610 & new_n5139;
  assign new_n12612 = ~new_n12589 & ~new_n12611;
  assign new_n12613 = ~new_n12612 & new_n5011;
  assign new_n12614 = ~new_n12567 & ~new_n12613;
  assign new_n12615 = ~new_n12614 & new_n5031;
  assign new_n12616 = ~new_n12521 & ~new_n12615;
  assign new_n12617 = ~new_n5077 & ~new_n12616;
  assign new_n12618 = ~new_n5207 & n2075;
  assign new_n12619 = n2107 & new_n5207;
  assign new_n12620 = ~new_n12618 & ~new_n12619;
  assign new_n12621 = ~new_n5243 & ~new_n12620;
  assign new_n12622 = ~new_n5207 & n2139;
  assign new_n12623 = n2171 & new_n5207;
  assign new_n12624 = ~new_n12622 & ~new_n12623;
  assign new_n12625 = ~new_n12624 & new_n5243;
  assign new_n12626 = ~new_n12621 & ~new_n12625;
  assign new_n12627 = ~new_n5170 & ~new_n12626;
  assign new_n12628 = ~new_n5207 & n2203;
  assign new_n12629 = n2235 & new_n5207;
  assign new_n12630 = ~new_n12628 & ~new_n12629;
  assign new_n12631 = ~new_n5243 & ~new_n12630;
  assign new_n12632 = ~new_n5207 & n2267;
  assign new_n12633 = n2299 & new_n5207;
  assign new_n12634 = ~new_n12632 & ~new_n12633;
  assign new_n12635 = ~new_n12634 & new_n5243;
  assign new_n12636 = ~new_n12631 & ~new_n12635;
  assign new_n12637 = ~new_n12636 & new_n5170;
  assign new_n12638 = ~new_n12627 & ~new_n12637;
  assign new_n12639 = ~new_n5139 & ~new_n12638;
  assign new_n12640 = ~new_n5207 & n2331;
  assign new_n12641 = n2363 & new_n5207;
  assign new_n12642 = ~new_n12640 & ~new_n12641;
  assign new_n12643 = ~new_n5243 & ~new_n12642;
  assign new_n12644 = ~new_n5207 & n2395;
  assign new_n12645 = n2427 & new_n5207;
  assign new_n12646 = ~new_n12644 & ~new_n12645;
  assign new_n12647 = ~new_n12646 & new_n5243;
  assign new_n12648 = ~new_n12643 & ~new_n12647;
  assign new_n12649 = ~new_n5170 & ~new_n12648;
  assign new_n12650 = ~new_n5207 & n2459;
  assign new_n12651 = n2491 & new_n5207;
  assign new_n12652 = ~new_n12650 & ~new_n12651;
  assign new_n12653 = ~new_n5243 & ~new_n12652;
  assign new_n12654 = ~new_n5207 & n2523;
  assign new_n12655 = n2555 & new_n5207;
  assign new_n12656 = ~new_n12654 & ~new_n12655;
  assign new_n12657 = ~new_n12656 & new_n5243;
  assign new_n12658 = ~new_n12653 & ~new_n12657;
  assign new_n12659 = ~new_n12658 & new_n5170;
  assign new_n12660 = ~new_n12649 & ~new_n12659;
  assign new_n12661 = ~new_n12660 & new_n5139;
  assign new_n12662 = ~new_n12639 & ~new_n12661;
  assign new_n12663 = ~new_n5011 & ~new_n12662;
  assign new_n12664 = ~new_n5207 & n2587;
  assign new_n12665 = n2619 & new_n5207;
  assign new_n12666 = ~new_n12664 & ~new_n12665;
  assign new_n12667 = ~new_n5243 & ~new_n12666;
  assign new_n12668 = ~new_n5207 & n2651;
  assign new_n12669 = n2683 & new_n5207;
  assign new_n12670 = ~new_n12668 & ~new_n12669;
  assign new_n12671 = ~new_n12670 & new_n5243;
  assign new_n12672 = ~new_n12667 & ~new_n12671;
  assign new_n12673 = ~new_n5170 & ~new_n12672;
  assign new_n12674 = ~new_n5207 & n2715;
  assign new_n12675 = n2747 & new_n5207;
  assign new_n12676 = ~new_n12674 & ~new_n12675;
  assign new_n12677 = ~new_n5243 & ~new_n12676;
  assign new_n12678 = ~new_n5207 & n2779;
  assign new_n12679 = n2811 & new_n5207;
  assign new_n12680 = ~new_n12678 & ~new_n12679;
  assign new_n12681 = ~new_n12680 & new_n5243;
  assign new_n12682 = ~new_n12677 & ~new_n12681;
  assign new_n12683 = ~new_n12682 & new_n5170;
  assign new_n12684 = ~new_n12673 & ~new_n12683;
  assign new_n12685 = ~new_n5139 & ~new_n12684;
  assign new_n12686 = ~new_n5207 & n2843;
  assign new_n12687 = n2875 & new_n5207;
  assign new_n12688 = ~new_n12686 & ~new_n12687;
  assign new_n12689 = ~new_n5243 & ~new_n12688;
  assign new_n12690 = ~new_n5207 & n2907;
  assign new_n12691 = n2939 & new_n5207;
  assign new_n12692 = ~new_n12690 & ~new_n12691;
  assign new_n12693 = ~new_n12692 & new_n5243;
  assign new_n12694 = ~new_n12689 & ~new_n12693;
  assign new_n12695 = ~new_n5170 & ~new_n12694;
  assign new_n12696 = ~new_n5207 & n2971;
  assign new_n12697 = n3003 & new_n5207;
  assign new_n12698 = ~new_n12696 & ~new_n12697;
  assign new_n12699 = ~new_n5243 & ~new_n12698;
  assign new_n12700 = ~new_n5207 & n3035;
  assign new_n12701 = n3067 & new_n5207;
  assign new_n12702 = ~new_n12700 & ~new_n12701;
  assign new_n12703 = ~new_n12702 & new_n5243;
  assign new_n12704 = ~new_n12699 & ~new_n12703;
  assign new_n12705 = ~new_n12704 & new_n5170;
  assign new_n12706 = ~new_n12695 & ~new_n12705;
  assign new_n12707 = ~new_n12706 & new_n5139;
  assign new_n12708 = ~new_n12685 & ~new_n12707;
  assign new_n12709 = ~new_n12708 & new_n5011;
  assign new_n12710 = ~new_n12663 & ~new_n12709;
  assign new_n12711 = ~new_n5031 & ~new_n12710;
  assign new_n12712 = ~new_n5207 & n3099;
  assign new_n12713 = n3131 & new_n5207;
  assign new_n12714 = ~new_n12712 & ~new_n12713;
  assign new_n12715 = ~new_n5243 & ~new_n12714;
  assign new_n12716 = ~new_n5207 & n3163;
  assign new_n12717 = n3195 & new_n5207;
  assign new_n12718 = ~new_n12716 & ~new_n12717;
  assign new_n12719 = ~new_n12718 & new_n5243;
  assign new_n12720 = ~new_n12715 & ~new_n12719;
  assign new_n12721 = ~new_n5170 & ~new_n12720;
  assign new_n12722 = ~new_n5207 & n3227;
  assign new_n12723 = n3259 & new_n5207;
  assign new_n12724 = ~new_n12722 & ~new_n12723;
  assign new_n12725 = ~new_n5243 & ~new_n12724;
  assign new_n12726 = ~new_n5207 & n3291;
  assign new_n12727 = n3323 & new_n5207;
  assign new_n12728 = ~new_n12726 & ~new_n12727;
  assign new_n12729 = ~new_n12728 & new_n5243;
  assign new_n12730 = ~new_n12725 & ~new_n12729;
  assign new_n12731 = ~new_n12730 & new_n5170;
  assign new_n12732 = ~new_n12721 & ~new_n12731;
  assign new_n12733 = ~new_n5139 & ~new_n12732;
  assign new_n12734 = ~new_n5207 & n3355;
  assign new_n12735 = n3387 & new_n5207;
  assign new_n12736 = ~new_n12734 & ~new_n12735;
  assign new_n12737 = ~new_n5243 & ~new_n12736;
  assign new_n12738 = ~new_n5207 & n3419;
  assign new_n12739 = n3451 & new_n5207;
  assign new_n12740 = ~new_n12738 & ~new_n12739;
  assign new_n12741 = ~new_n12740 & new_n5243;
  assign new_n12742 = ~new_n12737 & ~new_n12741;
  assign new_n12743 = ~new_n5170 & ~new_n12742;
  assign new_n12744 = ~new_n5207 & n3483;
  assign new_n12745 = n3515 & new_n5207;
  assign new_n12746 = ~new_n12744 & ~new_n12745;
  assign new_n12747 = ~new_n5243 & ~new_n12746;
  assign new_n12748 = ~new_n5207 & n3547;
  assign new_n12749 = n3579 & new_n5207;
  assign new_n12750 = ~new_n12748 & ~new_n12749;
  assign new_n12751 = ~new_n12750 & new_n5243;
  assign new_n12752 = ~new_n12747 & ~new_n12751;
  assign new_n12753 = ~new_n12752 & new_n5170;
  assign new_n12754 = ~new_n12743 & ~new_n12753;
  assign new_n12755 = ~new_n12754 & new_n5139;
  assign new_n12756 = ~new_n12733 & ~new_n12755;
  assign new_n12757 = ~new_n5011 & ~new_n12756;
  assign new_n12758 = ~new_n5207 & n3611;
  assign new_n12759 = n3643 & new_n5207;
  assign new_n12760 = ~new_n12758 & ~new_n12759;
  assign new_n12761 = ~new_n5243 & ~new_n12760;
  assign new_n12762 = ~new_n5207 & n3675;
  assign new_n12763 = n3707 & new_n5207;
  assign new_n12764 = ~new_n12762 & ~new_n12763;
  assign new_n12765 = ~new_n12764 & new_n5243;
  assign new_n12766 = ~new_n12761 & ~new_n12765;
  assign new_n12767 = ~new_n5170 & ~new_n12766;
  assign new_n12768 = ~new_n5207 & n3739;
  assign new_n12769 = n3771 & new_n5207;
  assign new_n12770 = ~new_n12768 & ~new_n12769;
  assign new_n12771 = ~new_n5243 & ~new_n12770;
  assign new_n12772 = ~new_n5207 & n3803;
  assign new_n12773 = n3835 & new_n5207;
  assign new_n12774 = ~new_n12772 & ~new_n12773;
  assign new_n12775 = ~new_n12774 & new_n5243;
  assign new_n12776 = ~new_n12771 & ~new_n12775;
  assign new_n12777 = ~new_n12776 & new_n5170;
  assign new_n12778 = ~new_n12767 & ~new_n12777;
  assign new_n12779 = ~new_n5139 & ~new_n12778;
  assign new_n12780 = ~new_n5207 & n3867;
  assign new_n12781 = n3899 & new_n5207;
  assign new_n12782 = ~new_n12780 & ~new_n12781;
  assign new_n12783 = ~new_n5243 & ~new_n12782;
  assign new_n12784 = ~new_n5207 & n3931;
  assign new_n12785 = n3963 & new_n5207;
  assign new_n12786 = ~new_n12784 & ~new_n12785;
  assign new_n12787 = ~new_n12786 & new_n5243;
  assign new_n12788 = ~new_n12783 & ~new_n12787;
  assign new_n12789 = ~new_n5170 & ~new_n12788;
  assign new_n12790 = ~new_n5207 & n3995;
  assign new_n12791 = n4027 & new_n5207;
  assign new_n12792 = ~new_n12790 & ~new_n12791;
  assign new_n12793 = ~new_n5243 & ~new_n12792;
  assign new_n12794 = ~new_n5207 & n4059;
  assign new_n12795 = n4091 & new_n5207;
  assign new_n12796 = ~new_n12794 & ~new_n12795;
  assign new_n12797 = ~new_n12796 & new_n5243;
  assign new_n12798 = ~new_n12793 & ~new_n12797;
  assign new_n12799 = ~new_n12798 & new_n5170;
  assign new_n12800 = ~new_n12789 & ~new_n12799;
  assign new_n12801 = ~new_n12800 & new_n5139;
  assign new_n12802 = ~new_n12779 & ~new_n12801;
  assign new_n12803 = ~new_n12802 & new_n5011;
  assign new_n12804 = ~new_n12757 & ~new_n12803;
  assign new_n12805 = ~new_n12804 & new_n5031;
  assign new_n12806 = ~new_n12711 & ~new_n12805;
  assign new_n12807 = ~new_n12806 & new_n5077;
  assign new_n12808 = ~new_n12617 & ~new_n12807;
  assign new_n12809 = ~new_n12808 & new_n8902;
  assign new_n12810 = ~new_n5207 & n2051;
  assign new_n12811 = n2083 & new_n5207;
  assign new_n12812 = ~new_n12810 & ~new_n12811;
  assign new_n12813 = ~new_n5243 & ~new_n12812;
  assign new_n12814 = ~new_n5207 & n2115;
  assign new_n12815 = n2147 & new_n5207;
  assign new_n12816 = ~new_n12814 & ~new_n12815;
  assign new_n12817 = ~new_n12816 & new_n5243;
  assign new_n12818 = ~new_n12813 & ~new_n12817;
  assign new_n12819 = ~new_n5170 & ~new_n12818;
  assign new_n12820 = ~new_n5207 & n2179;
  assign new_n12821 = n2211 & new_n5207;
  assign new_n12822 = ~new_n12820 & ~new_n12821;
  assign new_n12823 = ~new_n5243 & ~new_n12822;
  assign new_n12824 = ~new_n5207 & n2243;
  assign new_n12825 = n2275 & new_n5207;
  assign new_n12826 = ~new_n12824 & ~new_n12825;
  assign new_n12827 = ~new_n12826 & new_n5243;
  assign new_n12828 = ~new_n12823 & ~new_n12827;
  assign new_n12829 = ~new_n12828 & new_n5170;
  assign new_n12830 = ~new_n12819 & ~new_n12829;
  assign new_n12831 = ~new_n5139 & ~new_n12830;
  assign new_n12832 = ~new_n5207 & n2307;
  assign new_n12833 = n2339 & new_n5207;
  assign new_n12834 = ~new_n12832 & ~new_n12833;
  assign new_n12835 = ~new_n5243 & ~new_n12834;
  assign new_n12836 = ~new_n5207 & n2371;
  assign new_n12837 = n2403 & new_n5207;
  assign new_n12838 = ~new_n12836 & ~new_n12837;
  assign new_n12839 = ~new_n12838 & new_n5243;
  assign new_n12840 = ~new_n12835 & ~new_n12839;
  assign new_n12841 = ~new_n5170 & ~new_n12840;
  assign new_n12842 = ~new_n5207 & n2435;
  assign new_n12843 = n2467 & new_n5207;
  assign new_n12844 = ~new_n12842 & ~new_n12843;
  assign new_n12845 = ~new_n5243 & ~new_n12844;
  assign new_n12846 = ~new_n5207 & n2499;
  assign new_n12847 = n2531 & new_n5207;
  assign new_n12848 = ~new_n12846 & ~new_n12847;
  assign new_n12849 = ~new_n12848 & new_n5243;
  assign new_n12850 = ~new_n12845 & ~new_n12849;
  assign new_n12851 = ~new_n12850 & new_n5170;
  assign new_n12852 = ~new_n12841 & ~new_n12851;
  assign new_n12853 = ~new_n12852 & new_n5139;
  assign new_n12854 = ~new_n12831 & ~new_n12853;
  assign new_n12855 = ~new_n5011 & ~new_n12854;
  assign new_n12856 = ~new_n5207 & n2563;
  assign new_n12857 = n2595 & new_n5207;
  assign new_n12858 = ~new_n12856 & ~new_n12857;
  assign new_n12859 = ~new_n5243 & ~new_n12858;
  assign new_n12860 = ~new_n5207 & n2627;
  assign new_n12861 = n2659 & new_n5207;
  assign new_n12862 = ~new_n12860 & ~new_n12861;
  assign new_n12863 = ~new_n12862 & new_n5243;
  assign new_n12864 = ~new_n12859 & ~new_n12863;
  assign new_n12865 = ~new_n5170 & ~new_n12864;
  assign new_n12866 = ~new_n5207 & n2691;
  assign new_n12867 = n2723 & new_n5207;
  assign new_n12868 = ~new_n12866 & ~new_n12867;
  assign new_n12869 = ~new_n5243 & ~new_n12868;
  assign new_n12870 = ~new_n5207 & n2755;
  assign new_n12871 = n2787 & new_n5207;
  assign new_n12872 = ~new_n12870 & ~new_n12871;
  assign new_n12873 = ~new_n12872 & new_n5243;
  assign new_n12874 = ~new_n12869 & ~new_n12873;
  assign new_n12875 = ~new_n12874 & new_n5170;
  assign new_n12876 = ~new_n12865 & ~new_n12875;
  assign new_n12877 = ~new_n5139 & ~new_n12876;
  assign new_n12878 = ~new_n5207 & n2819;
  assign new_n12879 = n2851 & new_n5207;
  assign new_n12880 = ~new_n12878 & ~new_n12879;
  assign new_n12881 = ~new_n5243 & ~new_n12880;
  assign new_n12882 = ~new_n5207 & n2883;
  assign new_n12883 = n2915 & new_n5207;
  assign new_n12884 = ~new_n12882 & ~new_n12883;
  assign new_n12885 = ~new_n12884 & new_n5243;
  assign new_n12886 = ~new_n12881 & ~new_n12885;
  assign new_n12887 = ~new_n5170 & ~new_n12886;
  assign new_n12888 = ~new_n5207 & n2947;
  assign new_n12889 = n2979 & new_n5207;
  assign new_n12890 = ~new_n12888 & ~new_n12889;
  assign new_n12891 = ~new_n5243 & ~new_n12890;
  assign new_n12892 = ~new_n5207 & n3011;
  assign new_n12893 = n3043 & new_n5207;
  assign new_n12894 = ~new_n12892 & ~new_n12893;
  assign new_n12895 = ~new_n12894 & new_n5243;
  assign new_n12896 = ~new_n12891 & ~new_n12895;
  assign new_n12897 = ~new_n12896 & new_n5170;
  assign new_n12898 = ~new_n12887 & ~new_n12897;
  assign new_n12899 = ~new_n12898 & new_n5139;
  assign new_n12900 = ~new_n12877 & ~new_n12899;
  assign new_n12901 = ~new_n12900 & new_n5011;
  assign new_n12902 = ~new_n12855 & ~new_n12901;
  assign new_n12903 = ~new_n5031 & ~new_n12902;
  assign new_n12904 = ~new_n5207 & n3075;
  assign new_n12905 = n3107 & new_n5207;
  assign new_n12906 = ~new_n12904 & ~new_n12905;
  assign new_n12907 = ~new_n5243 & ~new_n12906;
  assign new_n12908 = ~new_n5207 & n3139;
  assign new_n12909 = n3171 & new_n5207;
  assign new_n12910 = ~new_n12908 & ~new_n12909;
  assign new_n12911 = ~new_n12910 & new_n5243;
  assign new_n12912 = ~new_n12907 & ~new_n12911;
  assign new_n12913 = ~new_n5170 & ~new_n12912;
  assign new_n12914 = ~new_n5207 & n3203;
  assign new_n12915 = n3235 & new_n5207;
  assign new_n12916 = ~new_n12914 & ~new_n12915;
  assign new_n12917 = ~new_n5243 & ~new_n12916;
  assign new_n12918 = ~new_n5207 & n3267;
  assign new_n12919 = n3299 & new_n5207;
  assign new_n12920 = ~new_n12918 & ~new_n12919;
  assign new_n12921 = ~new_n12920 & new_n5243;
  assign new_n12922 = ~new_n12917 & ~new_n12921;
  assign new_n12923 = ~new_n12922 & new_n5170;
  assign new_n12924 = ~new_n12913 & ~new_n12923;
  assign new_n12925 = ~new_n5139 & ~new_n12924;
  assign new_n12926 = ~new_n5207 & n3331;
  assign new_n12927 = n3363 & new_n5207;
  assign new_n12928 = ~new_n12926 & ~new_n12927;
  assign new_n12929 = ~new_n5243 & ~new_n12928;
  assign new_n12930 = ~new_n5207 & n3395;
  assign new_n12931 = n3427 & new_n5207;
  assign new_n12932 = ~new_n12930 & ~new_n12931;
  assign new_n12933 = ~new_n12932 & new_n5243;
  assign new_n12934 = ~new_n12929 & ~new_n12933;
  assign new_n12935 = ~new_n5170 & ~new_n12934;
  assign new_n12936 = ~new_n5207 & n3459;
  assign new_n12937 = n3491 & new_n5207;
  assign new_n12938 = ~new_n12936 & ~new_n12937;
  assign new_n12939 = ~new_n5243 & ~new_n12938;
  assign new_n12940 = ~new_n5207 & n3523;
  assign new_n12941 = n3555 & new_n5207;
  assign new_n12942 = ~new_n12940 & ~new_n12941;
  assign new_n12943 = ~new_n12942 & new_n5243;
  assign new_n12944 = ~new_n12939 & ~new_n12943;
  assign new_n12945 = ~new_n12944 & new_n5170;
  assign new_n12946 = ~new_n12935 & ~new_n12945;
  assign new_n12947 = ~new_n12946 & new_n5139;
  assign new_n12948 = ~new_n12925 & ~new_n12947;
  assign new_n12949 = ~new_n5011 & ~new_n12948;
  assign new_n12950 = ~new_n5207 & n3587;
  assign new_n12951 = n3619 & new_n5207;
  assign new_n12952 = ~new_n12950 & ~new_n12951;
  assign new_n12953 = ~new_n5243 & ~new_n12952;
  assign new_n12954 = ~new_n5207 & n3651;
  assign new_n12955 = n3683 & new_n5207;
  assign new_n12956 = ~new_n12954 & ~new_n12955;
  assign new_n12957 = ~new_n12956 & new_n5243;
  assign new_n12958 = ~new_n12953 & ~new_n12957;
  assign new_n12959 = ~new_n5170 & ~new_n12958;
  assign new_n12960 = ~new_n5207 & n3715;
  assign new_n12961 = n3747 & new_n5207;
  assign new_n12962 = ~new_n12960 & ~new_n12961;
  assign new_n12963 = ~new_n5243 & ~new_n12962;
  assign new_n12964 = ~new_n5207 & n3779;
  assign new_n12965 = n3811 & new_n5207;
  assign new_n12966 = ~new_n12964 & ~new_n12965;
  assign new_n12967 = ~new_n12966 & new_n5243;
  assign new_n12968 = ~new_n12963 & ~new_n12967;
  assign new_n12969 = ~new_n12968 & new_n5170;
  assign new_n12970 = ~new_n12959 & ~new_n12969;
  assign new_n12971 = ~new_n5139 & ~new_n12970;
  assign new_n12972 = ~new_n5207 & n3843;
  assign new_n12973 = n3875 & new_n5207;
  assign new_n12974 = ~new_n12972 & ~new_n12973;
  assign new_n12975 = ~new_n5243 & ~new_n12974;
  assign new_n12976 = ~new_n5207 & n3907;
  assign new_n12977 = n3939 & new_n5207;
  assign new_n12978 = ~new_n12976 & ~new_n12977;
  assign new_n12979 = ~new_n12978 & new_n5243;
  assign new_n12980 = ~new_n12975 & ~new_n12979;
  assign new_n12981 = ~new_n5170 & ~new_n12980;
  assign new_n12982 = ~new_n5207 & n3971;
  assign new_n12983 = n4003 & new_n5207;
  assign new_n12984 = ~new_n12982 & ~new_n12983;
  assign new_n12985 = ~new_n5243 & ~new_n12984;
  assign new_n12986 = ~new_n5207 & n4035;
  assign new_n12987 = n4067 & new_n5207;
  assign new_n12988 = ~new_n12986 & ~new_n12987;
  assign new_n12989 = ~new_n12988 & new_n5243;
  assign new_n12990 = ~new_n12985 & ~new_n12989;
  assign new_n12991 = ~new_n12990 & new_n5170;
  assign new_n12992 = ~new_n12981 & ~new_n12991;
  assign new_n12993 = ~new_n12992 & new_n5139;
  assign new_n12994 = ~new_n12971 & ~new_n12993;
  assign new_n12995 = ~new_n12994 & new_n5011;
  assign new_n12996 = ~new_n12949 & ~new_n12995;
  assign new_n12997 = ~new_n12996 & new_n5031;
  assign new_n12998 = ~new_n12903 & ~new_n12997;
  assign new_n12999 = ~new_n12998 & new_n5114;
  assign new_n13000 = ~new_n5462 & ~new_n12616;
  assign new_n13001 = ~new_n12999 & ~new_n13000;
  assign new_n13002 = ~new_n5207 & n2067;
  assign new_n13003 = n2099 & new_n5207;
  assign new_n13004 = ~new_n13002 & ~new_n13003;
  assign new_n13005 = ~new_n5243 & ~new_n13004;
  assign new_n13006 = ~new_n5207 & n2131;
  assign new_n13007 = n2163 & new_n5207;
  assign new_n13008 = ~new_n13006 & ~new_n13007;
  assign new_n13009 = ~new_n13008 & new_n5243;
  assign new_n13010 = ~new_n13005 & ~new_n13009;
  assign new_n13011 = ~new_n5170 & ~new_n13010;
  assign new_n13012 = ~new_n5207 & n2195;
  assign new_n13013 = n2227 & new_n5207;
  assign new_n13014 = ~new_n13012 & ~new_n13013;
  assign new_n13015 = ~new_n5243 & ~new_n13014;
  assign new_n13016 = ~new_n5207 & n2259;
  assign new_n13017 = n2291 & new_n5207;
  assign new_n13018 = ~new_n13016 & ~new_n13017;
  assign new_n13019 = ~new_n13018 & new_n5243;
  assign new_n13020 = ~new_n13015 & ~new_n13019;
  assign new_n13021 = ~new_n13020 & new_n5170;
  assign new_n13022 = ~new_n13011 & ~new_n13021;
  assign new_n13023 = ~new_n5139 & ~new_n13022;
  assign new_n13024 = ~new_n5207 & n2323;
  assign new_n13025 = n2355 & new_n5207;
  assign new_n13026 = ~new_n13024 & ~new_n13025;
  assign new_n13027 = ~new_n5243 & ~new_n13026;
  assign new_n13028 = ~new_n5207 & n2387;
  assign new_n13029 = n2419 & new_n5207;
  assign new_n13030 = ~new_n13028 & ~new_n13029;
  assign new_n13031 = ~new_n13030 & new_n5243;
  assign new_n13032 = ~new_n13027 & ~new_n13031;
  assign new_n13033 = ~new_n5170 & ~new_n13032;
  assign new_n13034 = ~new_n5207 & n2451;
  assign new_n13035 = n2483 & new_n5207;
  assign new_n13036 = ~new_n13034 & ~new_n13035;
  assign new_n13037 = ~new_n5243 & ~new_n13036;
  assign new_n13038 = ~new_n5207 & n2515;
  assign new_n13039 = n2547 & new_n5207;
  assign new_n13040 = ~new_n13038 & ~new_n13039;
  assign new_n13041 = ~new_n13040 & new_n5243;
  assign new_n13042 = ~new_n13037 & ~new_n13041;
  assign new_n13043 = ~new_n13042 & new_n5170;
  assign new_n13044 = ~new_n13033 & ~new_n13043;
  assign new_n13045 = ~new_n13044 & new_n5139;
  assign new_n13046 = ~new_n13023 & ~new_n13045;
  assign new_n13047 = ~new_n5011 & ~new_n13046;
  assign new_n13048 = ~new_n5207 & n2579;
  assign new_n13049 = n2611 & new_n5207;
  assign new_n13050 = ~new_n13048 & ~new_n13049;
  assign new_n13051 = ~new_n5243 & ~new_n13050;
  assign new_n13052 = ~new_n5207 & n2643;
  assign new_n13053 = n2675 & new_n5207;
  assign new_n13054 = ~new_n13052 & ~new_n13053;
  assign new_n13055 = ~new_n13054 & new_n5243;
  assign new_n13056 = ~new_n13051 & ~new_n13055;
  assign new_n13057 = ~new_n5170 & ~new_n13056;
  assign new_n13058 = ~new_n5207 & n2707;
  assign new_n13059 = n2739 & new_n5207;
  assign new_n13060 = ~new_n13058 & ~new_n13059;
  assign new_n13061 = ~new_n5243 & ~new_n13060;
  assign new_n13062 = ~new_n5207 & n2771;
  assign new_n13063 = n2803 & new_n5207;
  assign new_n13064 = ~new_n13062 & ~new_n13063;
  assign new_n13065 = ~new_n13064 & new_n5243;
  assign new_n13066 = ~new_n13061 & ~new_n13065;
  assign new_n13067 = ~new_n13066 & new_n5170;
  assign new_n13068 = ~new_n13057 & ~new_n13067;
  assign new_n13069 = ~new_n5139 & ~new_n13068;
  assign new_n13070 = ~new_n5207 & n2835;
  assign new_n13071 = n2867 & new_n5207;
  assign new_n13072 = ~new_n13070 & ~new_n13071;
  assign new_n13073 = ~new_n5243 & ~new_n13072;
  assign new_n13074 = ~new_n5207 & n2899;
  assign new_n13075 = n2931 & new_n5207;
  assign new_n13076 = ~new_n13074 & ~new_n13075;
  assign new_n13077 = ~new_n13076 & new_n5243;
  assign new_n13078 = ~new_n13073 & ~new_n13077;
  assign new_n13079 = ~new_n5170 & ~new_n13078;
  assign new_n13080 = ~new_n5207 & n2963;
  assign new_n13081 = n2995 & new_n5207;
  assign new_n13082 = ~new_n13080 & ~new_n13081;
  assign new_n13083 = ~new_n5243 & ~new_n13082;
  assign new_n13084 = ~new_n5207 & n3027;
  assign new_n13085 = n3059 & new_n5207;
  assign new_n13086 = ~new_n13084 & ~new_n13085;
  assign new_n13087 = ~new_n13086 & new_n5243;
  assign new_n13088 = ~new_n13083 & ~new_n13087;
  assign new_n13089 = ~new_n13088 & new_n5170;
  assign new_n13090 = ~new_n13079 & ~new_n13089;
  assign new_n13091 = ~new_n13090 & new_n5139;
  assign new_n13092 = ~new_n13069 & ~new_n13091;
  assign new_n13093 = ~new_n13092 & new_n5011;
  assign new_n13094 = ~new_n13047 & ~new_n13093;
  assign new_n13095 = ~new_n5031 & ~new_n13094;
  assign new_n13096 = ~new_n5207 & n3091;
  assign new_n13097 = n3123 & new_n5207;
  assign new_n13098 = ~new_n13096 & ~new_n13097;
  assign new_n13099 = ~new_n5243 & ~new_n13098;
  assign new_n13100 = ~new_n5207 & n3155;
  assign new_n13101 = n3187 & new_n5207;
  assign new_n13102 = ~new_n13100 & ~new_n13101;
  assign new_n13103 = ~new_n13102 & new_n5243;
  assign new_n13104 = ~new_n13099 & ~new_n13103;
  assign new_n13105 = ~new_n5170 & ~new_n13104;
  assign new_n13106 = ~new_n5207 & n3219;
  assign new_n13107 = n3251 & new_n5207;
  assign new_n13108 = ~new_n13106 & ~new_n13107;
  assign new_n13109 = ~new_n5243 & ~new_n13108;
  assign new_n13110 = ~new_n5207 & n3283;
  assign new_n13111 = n3315 & new_n5207;
  assign new_n13112 = ~new_n13110 & ~new_n13111;
  assign new_n13113 = ~new_n13112 & new_n5243;
  assign new_n13114 = ~new_n13109 & ~new_n13113;
  assign new_n13115 = ~new_n13114 & new_n5170;
  assign new_n13116 = ~new_n13105 & ~new_n13115;
  assign new_n13117 = ~new_n5139 & ~new_n13116;
  assign new_n13118 = ~new_n5207 & n3347;
  assign new_n13119 = n3379 & new_n5207;
  assign new_n13120 = ~new_n13118 & ~new_n13119;
  assign new_n13121 = ~new_n5243 & ~new_n13120;
  assign new_n13122 = ~new_n5207 & n3411;
  assign new_n13123 = n3443 & new_n5207;
  assign new_n13124 = ~new_n13122 & ~new_n13123;
  assign new_n13125 = ~new_n13124 & new_n5243;
  assign new_n13126 = ~new_n13121 & ~new_n13125;
  assign new_n13127 = ~new_n5170 & ~new_n13126;
  assign new_n13128 = ~new_n5207 & n3475;
  assign new_n13129 = n3507 & new_n5207;
  assign new_n13130 = ~new_n13128 & ~new_n13129;
  assign new_n13131 = ~new_n5243 & ~new_n13130;
  assign new_n13132 = ~new_n5207 & n3539;
  assign new_n13133 = n3571 & new_n5207;
  assign new_n13134 = ~new_n13132 & ~new_n13133;
  assign new_n13135 = ~new_n13134 & new_n5243;
  assign new_n13136 = ~new_n13131 & ~new_n13135;
  assign new_n13137 = ~new_n13136 & new_n5170;
  assign new_n13138 = ~new_n13127 & ~new_n13137;
  assign new_n13139 = ~new_n13138 & new_n5139;
  assign new_n13140 = ~new_n13117 & ~new_n13139;
  assign new_n13141 = ~new_n5011 & ~new_n13140;
  assign new_n13142 = ~new_n5207 & n3603;
  assign new_n13143 = n3635 & new_n5207;
  assign new_n13144 = ~new_n13142 & ~new_n13143;
  assign new_n13145 = ~new_n5243 & ~new_n13144;
  assign new_n13146 = ~new_n5207 & n3667;
  assign new_n13147 = n3699 & new_n5207;
  assign new_n13148 = ~new_n13146 & ~new_n13147;
  assign new_n13149 = ~new_n13148 & new_n5243;
  assign new_n13150 = ~new_n13145 & ~new_n13149;
  assign new_n13151 = ~new_n5170 & ~new_n13150;
  assign new_n13152 = ~new_n5207 & n3731;
  assign new_n13153 = n3763 & new_n5207;
  assign new_n13154 = ~new_n13152 & ~new_n13153;
  assign new_n13155 = ~new_n5243 & ~new_n13154;
  assign new_n13156 = ~new_n5207 & n3795;
  assign new_n13157 = n3827 & new_n5207;
  assign new_n13158 = ~new_n13156 & ~new_n13157;
  assign new_n13159 = ~new_n13158 & new_n5243;
  assign new_n13160 = ~new_n13155 & ~new_n13159;
  assign new_n13161 = ~new_n13160 & new_n5170;
  assign new_n13162 = ~new_n13151 & ~new_n13161;
  assign new_n13163 = ~new_n5139 & ~new_n13162;
  assign new_n13164 = ~new_n5207 & n3859;
  assign new_n13165 = n3891 & new_n5207;
  assign new_n13166 = ~new_n13164 & ~new_n13165;
  assign new_n13167 = ~new_n5243 & ~new_n13166;
  assign new_n13168 = ~new_n5207 & n3923;
  assign new_n13169 = n3955 & new_n5207;
  assign new_n13170 = ~new_n13168 & ~new_n13169;
  assign new_n13171 = ~new_n13170 & new_n5243;
  assign new_n13172 = ~new_n13167 & ~new_n13171;
  assign new_n13173 = ~new_n5170 & ~new_n13172;
  assign new_n13174 = ~new_n5207 & n3987;
  assign new_n13175 = n4019 & new_n5207;
  assign new_n13176 = ~new_n13174 & ~new_n13175;
  assign new_n13177 = ~new_n5243 & ~new_n13176;
  assign new_n13178 = ~new_n5207 & n4051;
  assign new_n13179 = n4083 & new_n5207;
  assign new_n13180 = ~new_n13178 & ~new_n13179;
  assign new_n13181 = ~new_n13180 & new_n5243;
  assign new_n13182 = ~new_n13177 & ~new_n13181;
  assign new_n13183 = ~new_n13182 & new_n5170;
  assign new_n13184 = ~new_n13173 & ~new_n13183;
  assign new_n13185 = ~new_n13184 & new_n5139;
  assign new_n13186 = ~new_n13163 & ~new_n13185;
  assign new_n13187 = ~new_n13186 & new_n5011;
  assign new_n13188 = ~new_n13141 & ~new_n13187;
  assign new_n13189 = ~new_n13188 & new_n5031;
  assign new_n13190 = ~new_n13095 & ~new_n13189;
  assign new_n13191 = ~new_n5115 & ~new_n13190;
  assign new_n13192 = ~new_n5116 & ~new_n12806;
  assign new_n13193 = ~new_n13191 & ~new_n13192;
  assign new_n13194 = new_n13001 & new_n13193;
  assign new_n13195 = ~new_n9289 & ~new_n13194;
  assign new_n13196 = ~new_n12809 & ~new_n13195;
  assign new_n13197 = ~new_n13194 & new_n8900;
  assign new_n13198 = ~new_n12808 & new_n8901;
  assign new_n13199 = ~new_n13197 & ~new_n13198;
  assign new_n13200 = ~new_n12806 & new_n4150;
  assign new_n13201 = ~new_n5139 & ~new_n9302;
  assign new_n13202 = ~new_n13200 & ~new_n13201;
  assign new_n13203 = new_n13199 & new_n13202;
  assign new_n13204 = new_n13196 & new_n13203;
  assign new_n13205 = ~new_n13204 & new_n8515;
  assign new_n13206 = ~new_n5207 & n2058;
  assign new_n13207 = n2090 & new_n5207;
  assign new_n13208 = ~new_n13206 & ~new_n13207;
  assign new_n13209 = ~new_n5243 & ~new_n13208;
  assign new_n13210 = ~new_n5207 & n2122;
  assign new_n13211 = n2154 & new_n5207;
  assign new_n13212 = ~new_n13210 & ~new_n13211;
  assign new_n13213 = ~new_n13212 & new_n5243;
  assign new_n13214 = ~new_n13209 & ~new_n13213;
  assign new_n13215 = ~new_n5170 & ~new_n13214;
  assign new_n13216 = ~new_n5207 & n2186;
  assign new_n13217 = n2218 & new_n5207;
  assign new_n13218 = ~new_n13216 & ~new_n13217;
  assign new_n13219 = ~new_n5243 & ~new_n13218;
  assign new_n13220 = ~new_n5207 & n2250;
  assign new_n13221 = n2282 & new_n5207;
  assign new_n13222 = ~new_n13220 & ~new_n13221;
  assign new_n13223 = ~new_n13222 & new_n5243;
  assign new_n13224 = ~new_n13219 & ~new_n13223;
  assign new_n13225 = ~new_n13224 & new_n5170;
  assign new_n13226 = ~new_n13215 & ~new_n13225;
  assign new_n13227 = ~new_n5139 & ~new_n13226;
  assign new_n13228 = ~new_n5207 & n2314;
  assign new_n13229 = n2346 & new_n5207;
  assign new_n13230 = ~new_n13228 & ~new_n13229;
  assign new_n13231 = ~new_n5243 & ~new_n13230;
  assign new_n13232 = ~new_n5207 & n2378;
  assign new_n13233 = n2410 & new_n5207;
  assign new_n13234 = ~new_n13232 & ~new_n13233;
  assign new_n13235 = ~new_n13234 & new_n5243;
  assign new_n13236 = ~new_n13231 & ~new_n13235;
  assign new_n13237 = ~new_n5170 & ~new_n13236;
  assign new_n13238 = ~new_n5207 & n2442;
  assign new_n13239 = n2474 & new_n5207;
  assign new_n13240 = ~new_n13238 & ~new_n13239;
  assign new_n13241 = ~new_n5243 & ~new_n13240;
  assign new_n13242 = ~new_n5207 & n2506;
  assign new_n13243 = n2538 & new_n5207;
  assign new_n13244 = ~new_n13242 & ~new_n13243;
  assign new_n13245 = ~new_n13244 & new_n5243;
  assign new_n13246 = ~new_n13241 & ~new_n13245;
  assign new_n13247 = ~new_n13246 & new_n5170;
  assign new_n13248 = ~new_n13237 & ~new_n13247;
  assign new_n13249 = ~new_n13248 & new_n5139;
  assign new_n13250 = ~new_n13227 & ~new_n13249;
  assign new_n13251 = ~new_n5011 & ~new_n13250;
  assign new_n13252 = ~new_n5207 & n2570;
  assign new_n13253 = n2602 & new_n5207;
  assign new_n13254 = ~new_n13252 & ~new_n13253;
  assign new_n13255 = ~new_n5243 & ~new_n13254;
  assign new_n13256 = ~new_n5207 & n2634;
  assign new_n13257 = n2666 & new_n5207;
  assign new_n13258 = ~new_n13256 & ~new_n13257;
  assign new_n13259 = ~new_n13258 & new_n5243;
  assign new_n13260 = ~new_n13255 & ~new_n13259;
  assign new_n13261 = ~new_n5170 & ~new_n13260;
  assign new_n13262 = ~new_n5207 & n2698;
  assign new_n13263 = n2730 & new_n5207;
  assign new_n13264 = ~new_n13262 & ~new_n13263;
  assign new_n13265 = ~new_n5243 & ~new_n13264;
  assign new_n13266 = ~new_n5207 & n2762;
  assign new_n13267 = n2794 & new_n5207;
  assign new_n13268 = ~new_n13266 & ~new_n13267;
  assign new_n13269 = ~new_n13268 & new_n5243;
  assign new_n13270 = ~new_n13265 & ~new_n13269;
  assign new_n13271 = ~new_n13270 & new_n5170;
  assign new_n13272 = ~new_n13261 & ~new_n13271;
  assign new_n13273 = ~new_n5139 & ~new_n13272;
  assign new_n13274 = ~new_n5207 & n2826;
  assign new_n13275 = n2858 & new_n5207;
  assign new_n13276 = ~new_n13274 & ~new_n13275;
  assign new_n13277 = ~new_n5243 & ~new_n13276;
  assign new_n13278 = ~new_n5207 & n2890;
  assign new_n13279 = n2922 & new_n5207;
  assign new_n13280 = ~new_n13278 & ~new_n13279;
  assign new_n13281 = ~new_n13280 & new_n5243;
  assign new_n13282 = ~new_n13277 & ~new_n13281;
  assign new_n13283 = ~new_n5170 & ~new_n13282;
  assign new_n13284 = ~new_n5207 & n2954;
  assign new_n13285 = n2986 & new_n5207;
  assign new_n13286 = ~new_n13284 & ~new_n13285;
  assign new_n13287 = ~new_n5243 & ~new_n13286;
  assign new_n13288 = ~new_n5207 & n3018;
  assign new_n13289 = n3050 & new_n5207;
  assign new_n13290 = ~new_n13288 & ~new_n13289;
  assign new_n13291 = ~new_n13290 & new_n5243;
  assign new_n13292 = ~new_n13287 & ~new_n13291;
  assign new_n13293 = ~new_n13292 & new_n5170;
  assign new_n13294 = ~new_n13283 & ~new_n13293;
  assign new_n13295 = ~new_n13294 & new_n5139;
  assign new_n13296 = ~new_n13273 & ~new_n13295;
  assign new_n13297 = ~new_n13296 & new_n5011;
  assign new_n13298 = ~new_n13251 & ~new_n13297;
  assign new_n13299 = ~new_n5031 & ~new_n13298;
  assign new_n13300 = ~new_n5207 & n3082;
  assign new_n13301 = n3114 & new_n5207;
  assign new_n13302 = ~new_n13300 & ~new_n13301;
  assign new_n13303 = ~new_n5243 & ~new_n13302;
  assign new_n13304 = ~new_n5207 & n3146;
  assign new_n13305 = n3178 & new_n5207;
  assign new_n13306 = ~new_n13304 & ~new_n13305;
  assign new_n13307 = ~new_n13306 & new_n5243;
  assign new_n13308 = ~new_n13303 & ~new_n13307;
  assign new_n13309 = ~new_n5170 & ~new_n13308;
  assign new_n13310 = ~new_n5207 & n3210;
  assign new_n13311 = n3242 & new_n5207;
  assign new_n13312 = ~new_n13310 & ~new_n13311;
  assign new_n13313 = ~new_n5243 & ~new_n13312;
  assign new_n13314 = ~new_n5207 & n3274;
  assign new_n13315 = n3306 & new_n5207;
  assign new_n13316 = ~new_n13314 & ~new_n13315;
  assign new_n13317 = ~new_n13316 & new_n5243;
  assign new_n13318 = ~new_n13313 & ~new_n13317;
  assign new_n13319 = ~new_n13318 & new_n5170;
  assign new_n13320 = ~new_n13309 & ~new_n13319;
  assign new_n13321 = ~new_n5139 & ~new_n13320;
  assign new_n13322 = ~new_n5207 & n3338;
  assign new_n13323 = n3370 & new_n5207;
  assign new_n13324 = ~new_n13322 & ~new_n13323;
  assign new_n13325 = ~new_n5243 & ~new_n13324;
  assign new_n13326 = ~new_n5207 & n3402;
  assign new_n13327 = n3434 & new_n5207;
  assign new_n13328 = ~new_n13326 & ~new_n13327;
  assign new_n13329 = ~new_n13328 & new_n5243;
  assign new_n13330 = ~new_n13325 & ~new_n13329;
  assign new_n13331 = ~new_n5170 & ~new_n13330;
  assign new_n13332 = ~new_n5207 & n3466;
  assign new_n13333 = n3498 & new_n5207;
  assign new_n13334 = ~new_n13332 & ~new_n13333;
  assign new_n13335 = ~new_n5243 & ~new_n13334;
  assign new_n13336 = ~new_n5207 & n3530;
  assign new_n13337 = n3562 & new_n5207;
  assign new_n13338 = ~new_n13336 & ~new_n13337;
  assign new_n13339 = ~new_n13338 & new_n5243;
  assign new_n13340 = ~new_n13335 & ~new_n13339;
  assign new_n13341 = ~new_n13340 & new_n5170;
  assign new_n13342 = ~new_n13331 & ~new_n13341;
  assign new_n13343 = ~new_n13342 & new_n5139;
  assign new_n13344 = ~new_n13321 & ~new_n13343;
  assign new_n13345 = ~new_n5011 & ~new_n13344;
  assign new_n13346 = ~new_n5207 & n3594;
  assign new_n13347 = n3626 & new_n5207;
  assign new_n13348 = ~new_n13346 & ~new_n13347;
  assign new_n13349 = ~new_n5243 & ~new_n13348;
  assign new_n13350 = ~new_n5207 & n3658;
  assign new_n13351 = n3690 & new_n5207;
  assign new_n13352 = ~new_n13350 & ~new_n13351;
  assign new_n13353 = ~new_n13352 & new_n5243;
  assign new_n13354 = ~new_n13349 & ~new_n13353;
  assign new_n13355 = ~new_n5170 & ~new_n13354;
  assign new_n13356 = ~new_n5207 & n3722;
  assign new_n13357 = n3754 & new_n5207;
  assign new_n13358 = ~new_n13356 & ~new_n13357;
  assign new_n13359 = ~new_n5243 & ~new_n13358;
  assign new_n13360 = ~new_n5207 & n3786;
  assign new_n13361 = n3818 & new_n5207;
  assign new_n13362 = ~new_n13360 & ~new_n13361;
  assign new_n13363 = ~new_n13362 & new_n5243;
  assign new_n13364 = ~new_n13359 & ~new_n13363;
  assign new_n13365 = ~new_n13364 & new_n5170;
  assign new_n13366 = ~new_n13355 & ~new_n13365;
  assign new_n13367 = ~new_n5139 & ~new_n13366;
  assign new_n13368 = ~new_n5207 & n3850;
  assign new_n13369 = n3882 & new_n5207;
  assign new_n13370 = ~new_n13368 & ~new_n13369;
  assign new_n13371 = ~new_n5243 & ~new_n13370;
  assign new_n13372 = ~new_n5207 & n3914;
  assign new_n13373 = n3946 & new_n5207;
  assign new_n13374 = ~new_n13372 & ~new_n13373;
  assign new_n13375 = ~new_n13374 & new_n5243;
  assign new_n13376 = ~new_n13371 & ~new_n13375;
  assign new_n13377 = ~new_n5170 & ~new_n13376;
  assign new_n13378 = ~new_n5207 & n3978;
  assign new_n13379 = n4010 & new_n5207;
  assign new_n13380 = ~new_n13378 & ~new_n13379;
  assign new_n13381 = ~new_n5243 & ~new_n13380;
  assign new_n13382 = ~new_n5207 & n4042;
  assign new_n13383 = n4074 & new_n5207;
  assign new_n13384 = ~new_n13382 & ~new_n13383;
  assign new_n13385 = ~new_n13384 & new_n5243;
  assign new_n13386 = ~new_n13381 & ~new_n13385;
  assign new_n13387 = ~new_n13386 & new_n5170;
  assign new_n13388 = ~new_n13377 & ~new_n13387;
  assign new_n13389 = ~new_n13388 & new_n5139;
  assign new_n13390 = ~new_n13367 & ~new_n13389;
  assign new_n13391 = ~new_n13390 & new_n5011;
  assign new_n13392 = ~new_n13345 & ~new_n13391;
  assign new_n13393 = ~new_n13392 & new_n5031;
  assign new_n13394 = ~new_n13299 & ~new_n13393;
  assign new_n13395 = ~new_n5077 & ~new_n13394;
  assign new_n13396 = ~new_n5207 & n2074;
  assign new_n13397 = n2106 & new_n5207;
  assign new_n13398 = ~new_n13396 & ~new_n13397;
  assign new_n13399 = ~new_n5243 & ~new_n13398;
  assign new_n13400 = ~new_n5207 & n2138;
  assign new_n13401 = n2170 & new_n5207;
  assign new_n13402 = ~new_n13400 & ~new_n13401;
  assign new_n13403 = ~new_n13402 & new_n5243;
  assign new_n13404 = ~new_n13399 & ~new_n13403;
  assign new_n13405 = ~new_n5170 & ~new_n13404;
  assign new_n13406 = ~new_n5207 & n2202;
  assign new_n13407 = n2234 & new_n5207;
  assign new_n13408 = ~new_n13406 & ~new_n13407;
  assign new_n13409 = ~new_n5243 & ~new_n13408;
  assign new_n13410 = ~new_n5207 & n2266;
  assign new_n13411 = n2298 & new_n5207;
  assign new_n13412 = ~new_n13410 & ~new_n13411;
  assign new_n13413 = ~new_n13412 & new_n5243;
  assign new_n13414 = ~new_n13409 & ~new_n13413;
  assign new_n13415 = ~new_n13414 & new_n5170;
  assign new_n13416 = ~new_n13405 & ~new_n13415;
  assign new_n13417 = ~new_n5139 & ~new_n13416;
  assign new_n13418 = ~new_n5207 & n2330;
  assign new_n13419 = n2362 & new_n5207;
  assign new_n13420 = ~new_n13418 & ~new_n13419;
  assign new_n13421 = ~new_n5243 & ~new_n13420;
  assign new_n13422 = ~new_n5207 & n2394;
  assign new_n13423 = n2426 & new_n5207;
  assign new_n13424 = ~new_n13422 & ~new_n13423;
  assign new_n13425 = ~new_n13424 & new_n5243;
  assign new_n13426 = ~new_n13421 & ~new_n13425;
  assign new_n13427 = ~new_n5170 & ~new_n13426;
  assign new_n13428 = ~new_n5207 & n2458;
  assign new_n13429 = n2490 & new_n5207;
  assign new_n13430 = ~new_n13428 & ~new_n13429;
  assign new_n13431 = ~new_n5243 & ~new_n13430;
  assign new_n13432 = ~new_n5207 & n2522;
  assign new_n13433 = n2554 & new_n5207;
  assign new_n13434 = ~new_n13432 & ~new_n13433;
  assign new_n13435 = ~new_n13434 & new_n5243;
  assign new_n13436 = ~new_n13431 & ~new_n13435;
  assign new_n13437 = ~new_n13436 & new_n5170;
  assign new_n13438 = ~new_n13427 & ~new_n13437;
  assign new_n13439 = ~new_n13438 & new_n5139;
  assign new_n13440 = ~new_n13417 & ~new_n13439;
  assign new_n13441 = ~new_n5011 & ~new_n13440;
  assign new_n13442 = ~new_n5207 & n2586;
  assign new_n13443 = n2618 & new_n5207;
  assign new_n13444 = ~new_n13442 & ~new_n13443;
  assign new_n13445 = ~new_n5243 & ~new_n13444;
  assign new_n13446 = ~new_n5207 & n2650;
  assign new_n13447 = n2682 & new_n5207;
  assign new_n13448 = ~new_n13446 & ~new_n13447;
  assign new_n13449 = ~new_n13448 & new_n5243;
  assign new_n13450 = ~new_n13445 & ~new_n13449;
  assign new_n13451 = ~new_n5170 & ~new_n13450;
  assign new_n13452 = ~new_n5207 & n2714;
  assign new_n13453 = n2746 & new_n5207;
  assign new_n13454 = ~new_n13452 & ~new_n13453;
  assign new_n13455 = ~new_n5243 & ~new_n13454;
  assign new_n13456 = ~new_n5207 & n2778;
  assign new_n13457 = n2810 & new_n5207;
  assign new_n13458 = ~new_n13456 & ~new_n13457;
  assign new_n13459 = ~new_n13458 & new_n5243;
  assign new_n13460 = ~new_n13455 & ~new_n13459;
  assign new_n13461 = ~new_n13460 & new_n5170;
  assign new_n13462 = ~new_n13451 & ~new_n13461;
  assign new_n13463 = ~new_n5139 & ~new_n13462;
  assign new_n13464 = ~new_n5207 & n2842;
  assign new_n13465 = n2874 & new_n5207;
  assign new_n13466 = ~new_n13464 & ~new_n13465;
  assign new_n13467 = ~new_n5243 & ~new_n13466;
  assign new_n13468 = ~new_n5207 & n2906;
  assign new_n13469 = n2938 & new_n5207;
  assign new_n13470 = ~new_n13468 & ~new_n13469;
  assign new_n13471 = ~new_n13470 & new_n5243;
  assign new_n13472 = ~new_n13467 & ~new_n13471;
  assign new_n13473 = ~new_n5170 & ~new_n13472;
  assign new_n13474 = ~new_n5207 & n2970;
  assign new_n13475 = n3002 & new_n5207;
  assign new_n13476 = ~new_n13474 & ~new_n13475;
  assign new_n13477 = ~new_n5243 & ~new_n13476;
  assign new_n13478 = ~new_n5207 & n3034;
  assign new_n13479 = n3066 & new_n5207;
  assign new_n13480 = ~new_n13478 & ~new_n13479;
  assign new_n13481 = ~new_n13480 & new_n5243;
  assign new_n13482 = ~new_n13477 & ~new_n13481;
  assign new_n13483 = ~new_n13482 & new_n5170;
  assign new_n13484 = ~new_n13473 & ~new_n13483;
  assign new_n13485 = ~new_n13484 & new_n5139;
  assign new_n13486 = ~new_n13463 & ~new_n13485;
  assign new_n13487 = ~new_n13486 & new_n5011;
  assign new_n13488 = ~new_n13441 & ~new_n13487;
  assign new_n13489 = ~new_n5031 & ~new_n13488;
  assign new_n13490 = ~new_n5207 & n3098;
  assign new_n13491 = n3130 & new_n5207;
  assign new_n13492 = ~new_n13490 & ~new_n13491;
  assign new_n13493 = ~new_n5243 & ~new_n13492;
  assign new_n13494 = ~new_n5207 & n3162;
  assign new_n13495 = n3194 & new_n5207;
  assign new_n13496 = ~new_n13494 & ~new_n13495;
  assign new_n13497 = ~new_n13496 & new_n5243;
  assign new_n13498 = ~new_n13493 & ~new_n13497;
  assign new_n13499 = ~new_n5170 & ~new_n13498;
  assign new_n13500 = ~new_n5207 & n3226;
  assign new_n13501 = n3258 & new_n5207;
  assign new_n13502 = ~new_n13500 & ~new_n13501;
  assign new_n13503 = ~new_n5243 & ~new_n13502;
  assign new_n13504 = ~new_n5207 & n3290;
  assign new_n13505 = n3322 & new_n5207;
  assign new_n13506 = ~new_n13504 & ~new_n13505;
  assign new_n13507 = ~new_n13506 & new_n5243;
  assign new_n13508 = ~new_n13503 & ~new_n13507;
  assign new_n13509 = ~new_n13508 & new_n5170;
  assign new_n13510 = ~new_n13499 & ~new_n13509;
  assign new_n13511 = ~new_n5139 & ~new_n13510;
  assign new_n13512 = ~new_n5207 & n3354;
  assign new_n13513 = n3386 & new_n5207;
  assign new_n13514 = ~new_n13512 & ~new_n13513;
  assign new_n13515 = ~new_n5243 & ~new_n13514;
  assign new_n13516 = ~new_n5207 & n3418;
  assign new_n13517 = n3450 & new_n5207;
  assign new_n13518 = ~new_n13516 & ~new_n13517;
  assign new_n13519 = ~new_n13518 & new_n5243;
  assign new_n13520 = ~new_n13515 & ~new_n13519;
  assign new_n13521 = ~new_n5170 & ~new_n13520;
  assign new_n13522 = ~new_n5207 & n3482;
  assign new_n13523 = n3514 & new_n5207;
  assign new_n13524 = ~new_n13522 & ~new_n13523;
  assign new_n13525 = ~new_n5243 & ~new_n13524;
  assign new_n13526 = ~new_n5207 & n3546;
  assign new_n13527 = n3578 & new_n5207;
  assign new_n13528 = ~new_n13526 & ~new_n13527;
  assign new_n13529 = ~new_n13528 & new_n5243;
  assign new_n13530 = ~new_n13525 & ~new_n13529;
  assign new_n13531 = ~new_n13530 & new_n5170;
  assign new_n13532 = ~new_n13521 & ~new_n13531;
  assign new_n13533 = ~new_n13532 & new_n5139;
  assign new_n13534 = ~new_n13511 & ~new_n13533;
  assign new_n13535 = ~new_n5011 & ~new_n13534;
  assign new_n13536 = ~new_n5207 & n3610;
  assign new_n13537 = n3642 & new_n5207;
  assign new_n13538 = ~new_n13536 & ~new_n13537;
  assign new_n13539 = ~new_n5243 & ~new_n13538;
  assign new_n13540 = ~new_n5207 & n3674;
  assign new_n13541 = n3706 & new_n5207;
  assign new_n13542 = ~new_n13540 & ~new_n13541;
  assign new_n13543 = ~new_n13542 & new_n5243;
  assign new_n13544 = ~new_n13539 & ~new_n13543;
  assign new_n13545 = ~new_n5170 & ~new_n13544;
  assign new_n13546 = ~new_n5207 & n3738;
  assign new_n13547 = n3770 & new_n5207;
  assign new_n13548 = ~new_n13546 & ~new_n13547;
  assign new_n13549 = ~new_n5243 & ~new_n13548;
  assign new_n13550 = ~new_n5207 & n3802;
  assign new_n13551 = n3834 & new_n5207;
  assign new_n13552 = ~new_n13550 & ~new_n13551;
  assign new_n13553 = ~new_n13552 & new_n5243;
  assign new_n13554 = ~new_n13549 & ~new_n13553;
  assign new_n13555 = ~new_n13554 & new_n5170;
  assign new_n13556 = ~new_n13545 & ~new_n13555;
  assign new_n13557 = ~new_n5139 & ~new_n13556;
  assign new_n13558 = ~new_n5207 & n3866;
  assign new_n13559 = n3898 & new_n5207;
  assign new_n13560 = ~new_n13558 & ~new_n13559;
  assign new_n13561 = ~new_n5243 & ~new_n13560;
  assign new_n13562 = ~new_n5207 & n3930;
  assign new_n13563 = n3962 & new_n5207;
  assign new_n13564 = ~new_n13562 & ~new_n13563;
  assign new_n13565 = ~new_n13564 & new_n5243;
  assign new_n13566 = ~new_n13561 & ~new_n13565;
  assign new_n13567 = ~new_n5170 & ~new_n13566;
  assign new_n13568 = ~new_n5207 & n3994;
  assign new_n13569 = n4026 & new_n5207;
  assign new_n13570 = ~new_n13568 & ~new_n13569;
  assign new_n13571 = ~new_n5243 & ~new_n13570;
  assign new_n13572 = ~new_n5207 & n4058;
  assign new_n13573 = n4090 & new_n5207;
  assign new_n13574 = ~new_n13572 & ~new_n13573;
  assign new_n13575 = ~new_n13574 & new_n5243;
  assign new_n13576 = ~new_n13571 & ~new_n13575;
  assign new_n13577 = ~new_n13576 & new_n5170;
  assign new_n13578 = ~new_n13567 & ~new_n13577;
  assign new_n13579 = ~new_n13578 & new_n5139;
  assign new_n13580 = ~new_n13557 & ~new_n13579;
  assign new_n13581 = ~new_n13580 & new_n5011;
  assign new_n13582 = ~new_n13535 & ~new_n13581;
  assign new_n13583 = ~new_n13582 & new_n5031;
  assign new_n13584 = ~new_n13489 & ~new_n13583;
  assign new_n13585 = ~new_n13584 & new_n5077;
  assign new_n13586 = ~new_n13395 & ~new_n13585;
  assign new_n13587 = ~new_n13586 & new_n8902;
  assign new_n13588 = ~new_n5207 & n2050;
  assign new_n13589 = n2082 & new_n5207;
  assign new_n13590 = ~new_n13588 & ~new_n13589;
  assign new_n13591 = ~new_n5243 & ~new_n13590;
  assign new_n13592 = ~new_n5207 & n2114;
  assign new_n13593 = n2146 & new_n5207;
  assign new_n13594 = ~new_n13592 & ~new_n13593;
  assign new_n13595 = ~new_n13594 & new_n5243;
  assign new_n13596 = ~new_n13591 & ~new_n13595;
  assign new_n13597 = ~new_n5170 & ~new_n13596;
  assign new_n13598 = ~new_n5207 & n2178;
  assign new_n13599 = n2210 & new_n5207;
  assign new_n13600 = ~new_n13598 & ~new_n13599;
  assign new_n13601 = ~new_n5243 & ~new_n13600;
  assign new_n13602 = ~new_n5207 & n2242;
  assign new_n13603 = n2274 & new_n5207;
  assign new_n13604 = ~new_n13602 & ~new_n13603;
  assign new_n13605 = ~new_n13604 & new_n5243;
  assign new_n13606 = ~new_n13601 & ~new_n13605;
  assign new_n13607 = ~new_n13606 & new_n5170;
  assign new_n13608 = ~new_n13597 & ~new_n13607;
  assign new_n13609 = ~new_n5139 & ~new_n13608;
  assign new_n13610 = ~new_n5207 & n2306;
  assign new_n13611 = n2338 & new_n5207;
  assign new_n13612 = ~new_n13610 & ~new_n13611;
  assign new_n13613 = ~new_n5243 & ~new_n13612;
  assign new_n13614 = ~new_n5207 & n2370;
  assign new_n13615 = n2402 & new_n5207;
  assign new_n13616 = ~new_n13614 & ~new_n13615;
  assign new_n13617 = ~new_n13616 & new_n5243;
  assign new_n13618 = ~new_n13613 & ~new_n13617;
  assign new_n13619 = ~new_n5170 & ~new_n13618;
  assign new_n13620 = ~new_n5207 & n2434;
  assign new_n13621 = n2466 & new_n5207;
  assign new_n13622 = ~new_n13620 & ~new_n13621;
  assign new_n13623 = ~new_n5243 & ~new_n13622;
  assign new_n13624 = ~new_n5207 & n2498;
  assign new_n13625 = n2530 & new_n5207;
  assign new_n13626 = ~new_n13624 & ~new_n13625;
  assign new_n13627 = ~new_n13626 & new_n5243;
  assign new_n13628 = ~new_n13623 & ~new_n13627;
  assign new_n13629 = ~new_n13628 & new_n5170;
  assign new_n13630 = ~new_n13619 & ~new_n13629;
  assign new_n13631 = ~new_n13630 & new_n5139;
  assign new_n13632 = ~new_n13609 & ~new_n13631;
  assign new_n13633 = ~new_n5011 & ~new_n13632;
  assign new_n13634 = ~new_n5207 & n2562;
  assign new_n13635 = n2594 & new_n5207;
  assign new_n13636 = ~new_n13634 & ~new_n13635;
  assign new_n13637 = ~new_n5243 & ~new_n13636;
  assign new_n13638 = ~new_n5207 & n2626;
  assign new_n13639 = n2658 & new_n5207;
  assign new_n13640 = ~new_n13638 & ~new_n13639;
  assign new_n13641 = ~new_n13640 & new_n5243;
  assign new_n13642 = ~new_n13637 & ~new_n13641;
  assign new_n13643 = ~new_n5170 & ~new_n13642;
  assign new_n13644 = ~new_n5207 & n2690;
  assign new_n13645 = n2722 & new_n5207;
  assign new_n13646 = ~new_n13644 & ~new_n13645;
  assign new_n13647 = ~new_n5243 & ~new_n13646;
  assign new_n13648 = ~new_n5207 & n2754;
  assign new_n13649 = n2786 & new_n5207;
  assign new_n13650 = ~new_n13648 & ~new_n13649;
  assign new_n13651 = ~new_n13650 & new_n5243;
  assign new_n13652 = ~new_n13647 & ~new_n13651;
  assign new_n13653 = ~new_n13652 & new_n5170;
  assign new_n13654 = ~new_n13643 & ~new_n13653;
  assign new_n13655 = ~new_n5139 & ~new_n13654;
  assign new_n13656 = ~new_n5207 & n2818;
  assign new_n13657 = n2850 & new_n5207;
  assign new_n13658 = ~new_n13656 & ~new_n13657;
  assign new_n13659 = ~new_n5243 & ~new_n13658;
  assign new_n13660 = ~new_n5207 & n2882;
  assign new_n13661 = n2914 & new_n5207;
  assign new_n13662 = ~new_n13660 & ~new_n13661;
  assign new_n13663 = ~new_n13662 & new_n5243;
  assign new_n13664 = ~new_n13659 & ~new_n13663;
  assign new_n13665 = ~new_n5170 & ~new_n13664;
  assign new_n13666 = ~new_n5207 & n2946;
  assign new_n13667 = n2978 & new_n5207;
  assign new_n13668 = ~new_n13666 & ~new_n13667;
  assign new_n13669 = ~new_n5243 & ~new_n13668;
  assign new_n13670 = ~new_n5207 & n3010;
  assign new_n13671 = n3042 & new_n5207;
  assign new_n13672 = ~new_n13670 & ~new_n13671;
  assign new_n13673 = ~new_n13672 & new_n5243;
  assign new_n13674 = ~new_n13669 & ~new_n13673;
  assign new_n13675 = ~new_n13674 & new_n5170;
  assign new_n13676 = ~new_n13665 & ~new_n13675;
  assign new_n13677 = ~new_n13676 & new_n5139;
  assign new_n13678 = ~new_n13655 & ~new_n13677;
  assign new_n13679 = ~new_n13678 & new_n5011;
  assign new_n13680 = ~new_n13633 & ~new_n13679;
  assign new_n13681 = ~new_n5031 & ~new_n13680;
  assign new_n13682 = ~new_n5207 & n3074;
  assign new_n13683 = n3106 & new_n5207;
  assign new_n13684 = ~new_n13682 & ~new_n13683;
  assign new_n13685 = ~new_n5243 & ~new_n13684;
  assign new_n13686 = ~new_n5207 & n3138;
  assign new_n13687 = n3170 & new_n5207;
  assign new_n13688 = ~new_n13686 & ~new_n13687;
  assign new_n13689 = ~new_n13688 & new_n5243;
  assign new_n13690 = ~new_n13685 & ~new_n13689;
  assign new_n13691 = ~new_n5170 & ~new_n13690;
  assign new_n13692 = ~new_n5207 & n3202;
  assign new_n13693 = n3234 & new_n5207;
  assign new_n13694 = ~new_n13692 & ~new_n13693;
  assign new_n13695 = ~new_n5243 & ~new_n13694;
  assign new_n13696 = ~new_n5207 & n3266;
  assign new_n13697 = n3298 & new_n5207;
  assign new_n13698 = ~new_n13696 & ~new_n13697;
  assign new_n13699 = ~new_n13698 & new_n5243;
  assign new_n13700 = ~new_n13695 & ~new_n13699;
  assign new_n13701 = ~new_n13700 & new_n5170;
  assign new_n13702 = ~new_n13691 & ~new_n13701;
  assign new_n13703 = ~new_n5139 & ~new_n13702;
  assign new_n13704 = ~new_n5207 & n3330;
  assign new_n13705 = n3362 & new_n5207;
  assign new_n13706 = ~new_n13704 & ~new_n13705;
  assign new_n13707 = ~new_n5243 & ~new_n13706;
  assign new_n13708 = ~new_n5207 & n3394;
  assign new_n13709 = n3426 & new_n5207;
  assign new_n13710 = ~new_n13708 & ~new_n13709;
  assign new_n13711 = ~new_n13710 & new_n5243;
  assign new_n13712 = ~new_n13707 & ~new_n13711;
  assign new_n13713 = ~new_n5170 & ~new_n13712;
  assign new_n13714 = ~new_n5207 & n3458;
  assign new_n13715 = n3490 & new_n5207;
  assign new_n13716 = ~new_n13714 & ~new_n13715;
  assign new_n13717 = ~new_n5243 & ~new_n13716;
  assign new_n13718 = ~new_n5207 & n3522;
  assign new_n13719 = n3554 & new_n5207;
  assign new_n13720 = ~new_n13718 & ~new_n13719;
  assign new_n13721 = ~new_n13720 & new_n5243;
  assign new_n13722 = ~new_n13717 & ~new_n13721;
  assign new_n13723 = ~new_n13722 & new_n5170;
  assign new_n13724 = ~new_n13713 & ~new_n13723;
  assign new_n13725 = ~new_n13724 & new_n5139;
  assign new_n13726 = ~new_n13703 & ~new_n13725;
  assign new_n13727 = ~new_n5011 & ~new_n13726;
  assign new_n13728 = ~new_n5207 & n3586;
  assign new_n13729 = n3618 & new_n5207;
  assign new_n13730 = ~new_n13728 & ~new_n13729;
  assign new_n13731 = ~new_n5243 & ~new_n13730;
  assign new_n13732 = ~new_n5207 & n3650;
  assign new_n13733 = n3682 & new_n5207;
  assign new_n13734 = ~new_n13732 & ~new_n13733;
  assign new_n13735 = ~new_n13734 & new_n5243;
  assign new_n13736 = ~new_n13731 & ~new_n13735;
  assign new_n13737 = ~new_n5170 & ~new_n13736;
  assign new_n13738 = ~new_n5207 & n3714;
  assign new_n13739 = n3746 & new_n5207;
  assign new_n13740 = ~new_n13738 & ~new_n13739;
  assign new_n13741 = ~new_n5243 & ~new_n13740;
  assign new_n13742 = ~new_n5207 & n3778;
  assign new_n13743 = n3810 & new_n5207;
  assign new_n13744 = ~new_n13742 & ~new_n13743;
  assign new_n13745 = ~new_n13744 & new_n5243;
  assign new_n13746 = ~new_n13741 & ~new_n13745;
  assign new_n13747 = ~new_n13746 & new_n5170;
  assign new_n13748 = ~new_n13737 & ~new_n13747;
  assign new_n13749 = ~new_n5139 & ~new_n13748;
  assign new_n13750 = ~new_n5207 & n3842;
  assign new_n13751 = n3874 & new_n5207;
  assign new_n13752 = ~new_n13750 & ~new_n13751;
  assign new_n13753 = ~new_n5243 & ~new_n13752;
  assign new_n13754 = ~new_n5207 & n3906;
  assign new_n13755 = n3938 & new_n5207;
  assign new_n13756 = ~new_n13754 & ~new_n13755;
  assign new_n13757 = ~new_n13756 & new_n5243;
  assign new_n13758 = ~new_n13753 & ~new_n13757;
  assign new_n13759 = ~new_n5170 & ~new_n13758;
  assign new_n13760 = ~new_n5207 & n3970;
  assign new_n13761 = n4002 & new_n5207;
  assign new_n13762 = ~new_n13760 & ~new_n13761;
  assign new_n13763 = ~new_n5243 & ~new_n13762;
  assign new_n13764 = ~new_n5207 & n4034;
  assign new_n13765 = n4066 & new_n5207;
  assign new_n13766 = ~new_n13764 & ~new_n13765;
  assign new_n13767 = ~new_n13766 & new_n5243;
  assign new_n13768 = ~new_n13763 & ~new_n13767;
  assign new_n13769 = ~new_n13768 & new_n5170;
  assign new_n13770 = ~new_n13759 & ~new_n13769;
  assign new_n13771 = ~new_n13770 & new_n5139;
  assign new_n13772 = ~new_n13749 & ~new_n13771;
  assign new_n13773 = ~new_n13772 & new_n5011;
  assign new_n13774 = ~new_n13727 & ~new_n13773;
  assign new_n13775 = ~new_n13774 & new_n5031;
  assign new_n13776 = ~new_n13681 & ~new_n13775;
  assign new_n13777 = ~new_n13776 & new_n5114;
  assign new_n13778 = ~new_n5462 & ~new_n13394;
  assign new_n13779 = ~new_n13777 & ~new_n13778;
  assign new_n13780 = ~new_n5207 & n2066;
  assign new_n13781 = n2098 & new_n5207;
  assign new_n13782 = ~new_n13780 & ~new_n13781;
  assign new_n13783 = ~new_n5243 & ~new_n13782;
  assign new_n13784 = ~new_n5207 & n2130;
  assign new_n13785 = n2162 & new_n5207;
  assign new_n13786 = ~new_n13784 & ~new_n13785;
  assign new_n13787 = ~new_n13786 & new_n5243;
  assign new_n13788 = ~new_n13783 & ~new_n13787;
  assign new_n13789 = ~new_n5170 & ~new_n13788;
  assign new_n13790 = ~new_n5207 & n2194;
  assign new_n13791 = n2226 & new_n5207;
  assign new_n13792 = ~new_n13790 & ~new_n13791;
  assign new_n13793 = ~new_n5243 & ~new_n13792;
  assign new_n13794 = ~new_n5207 & n2258;
  assign new_n13795 = n2290 & new_n5207;
  assign new_n13796 = ~new_n13794 & ~new_n13795;
  assign new_n13797 = ~new_n13796 & new_n5243;
  assign new_n13798 = ~new_n13793 & ~new_n13797;
  assign new_n13799 = ~new_n13798 & new_n5170;
  assign new_n13800 = ~new_n13789 & ~new_n13799;
  assign new_n13801 = ~new_n5139 & ~new_n13800;
  assign new_n13802 = ~new_n5207 & n2322;
  assign new_n13803 = n2354 & new_n5207;
  assign new_n13804 = ~new_n13802 & ~new_n13803;
  assign new_n13805 = ~new_n5243 & ~new_n13804;
  assign new_n13806 = ~new_n5207 & n2386;
  assign new_n13807 = n2418 & new_n5207;
  assign new_n13808 = ~new_n13806 & ~new_n13807;
  assign new_n13809 = ~new_n13808 & new_n5243;
  assign new_n13810 = ~new_n13805 & ~new_n13809;
  assign new_n13811 = ~new_n5170 & ~new_n13810;
  assign new_n13812 = ~new_n5207 & n2450;
  assign new_n13813 = n2482 & new_n5207;
  assign new_n13814 = ~new_n13812 & ~new_n13813;
  assign new_n13815 = ~new_n5243 & ~new_n13814;
  assign new_n13816 = ~new_n5207 & n2514;
  assign new_n13817 = n2546 & new_n5207;
  assign new_n13818 = ~new_n13816 & ~new_n13817;
  assign new_n13819 = ~new_n13818 & new_n5243;
  assign new_n13820 = ~new_n13815 & ~new_n13819;
  assign new_n13821 = ~new_n13820 & new_n5170;
  assign new_n13822 = ~new_n13811 & ~new_n13821;
  assign new_n13823 = ~new_n13822 & new_n5139;
  assign new_n13824 = ~new_n13801 & ~new_n13823;
  assign new_n13825 = ~new_n5011 & ~new_n13824;
  assign new_n13826 = ~new_n5207 & n2578;
  assign new_n13827 = n2610 & new_n5207;
  assign new_n13828 = ~new_n13826 & ~new_n13827;
  assign new_n13829 = ~new_n5243 & ~new_n13828;
  assign new_n13830 = ~new_n5207 & n2642;
  assign new_n13831 = n2674 & new_n5207;
  assign new_n13832 = ~new_n13830 & ~new_n13831;
  assign new_n13833 = ~new_n13832 & new_n5243;
  assign new_n13834 = ~new_n13829 & ~new_n13833;
  assign new_n13835 = ~new_n5170 & ~new_n13834;
  assign new_n13836 = ~new_n5207 & n2706;
  assign new_n13837 = n2738 & new_n5207;
  assign new_n13838 = ~new_n13836 & ~new_n13837;
  assign new_n13839 = ~new_n5243 & ~new_n13838;
  assign new_n13840 = ~new_n5207 & n2770;
  assign new_n13841 = n2802 & new_n5207;
  assign new_n13842 = ~new_n13840 & ~new_n13841;
  assign new_n13843 = ~new_n13842 & new_n5243;
  assign new_n13844 = ~new_n13839 & ~new_n13843;
  assign new_n13845 = ~new_n13844 & new_n5170;
  assign new_n13846 = ~new_n13835 & ~new_n13845;
  assign new_n13847 = ~new_n5139 & ~new_n13846;
  assign new_n13848 = ~new_n5207 & n2834;
  assign new_n13849 = n2866 & new_n5207;
  assign new_n13850 = ~new_n13848 & ~new_n13849;
  assign new_n13851 = ~new_n5243 & ~new_n13850;
  assign new_n13852 = ~new_n5207 & n2898;
  assign new_n13853 = n2930 & new_n5207;
  assign new_n13854 = ~new_n13852 & ~new_n13853;
  assign new_n13855 = ~new_n13854 & new_n5243;
  assign new_n13856 = ~new_n13851 & ~new_n13855;
  assign new_n13857 = ~new_n5170 & ~new_n13856;
  assign new_n13858 = ~new_n5207 & n2962;
  assign new_n13859 = n2994 & new_n5207;
  assign new_n13860 = ~new_n13858 & ~new_n13859;
  assign new_n13861 = ~new_n5243 & ~new_n13860;
  assign new_n13862 = ~new_n5207 & n3026;
  assign new_n13863 = n3058 & new_n5207;
  assign new_n13864 = ~new_n13862 & ~new_n13863;
  assign new_n13865 = ~new_n13864 & new_n5243;
  assign new_n13866 = ~new_n13861 & ~new_n13865;
  assign new_n13867 = ~new_n13866 & new_n5170;
  assign new_n13868 = ~new_n13857 & ~new_n13867;
  assign new_n13869 = ~new_n13868 & new_n5139;
  assign new_n13870 = ~new_n13847 & ~new_n13869;
  assign new_n13871 = ~new_n13870 & new_n5011;
  assign new_n13872 = ~new_n13825 & ~new_n13871;
  assign new_n13873 = ~new_n5031 & ~new_n13872;
  assign new_n13874 = ~new_n5207 & n3090;
  assign new_n13875 = n3122 & new_n5207;
  assign new_n13876 = ~new_n13874 & ~new_n13875;
  assign new_n13877 = ~new_n5243 & ~new_n13876;
  assign new_n13878 = ~new_n5207 & n3154;
  assign new_n13879 = n3186 & new_n5207;
  assign new_n13880 = ~new_n13878 & ~new_n13879;
  assign new_n13881 = ~new_n13880 & new_n5243;
  assign new_n13882 = ~new_n13877 & ~new_n13881;
  assign new_n13883 = ~new_n5170 & ~new_n13882;
  assign new_n13884 = ~new_n5207 & n3218;
  assign new_n13885 = n3250 & new_n5207;
  assign new_n13886 = ~new_n13884 & ~new_n13885;
  assign new_n13887 = ~new_n5243 & ~new_n13886;
  assign new_n13888 = ~new_n5207 & n3282;
  assign new_n13889 = n3314 & new_n5207;
  assign new_n13890 = ~new_n13888 & ~new_n13889;
  assign new_n13891 = ~new_n13890 & new_n5243;
  assign new_n13892 = ~new_n13887 & ~new_n13891;
  assign new_n13893 = ~new_n13892 & new_n5170;
  assign new_n13894 = ~new_n13883 & ~new_n13893;
  assign new_n13895 = ~new_n5139 & ~new_n13894;
  assign new_n13896 = ~new_n5207 & n3346;
  assign new_n13897 = n3378 & new_n5207;
  assign new_n13898 = ~new_n13896 & ~new_n13897;
  assign new_n13899 = ~new_n5243 & ~new_n13898;
  assign new_n13900 = ~new_n5207 & n3410;
  assign new_n13901 = n3442 & new_n5207;
  assign new_n13902 = ~new_n13900 & ~new_n13901;
  assign new_n13903 = ~new_n13902 & new_n5243;
  assign new_n13904 = ~new_n13899 & ~new_n13903;
  assign new_n13905 = ~new_n5170 & ~new_n13904;
  assign new_n13906 = ~new_n5207 & n3474;
  assign new_n13907 = n3506 & new_n5207;
  assign new_n13908 = ~new_n13906 & ~new_n13907;
  assign new_n13909 = ~new_n5243 & ~new_n13908;
  assign new_n13910 = ~new_n5207 & n3538;
  assign new_n13911 = n3570 & new_n5207;
  assign new_n13912 = ~new_n13910 & ~new_n13911;
  assign new_n13913 = ~new_n13912 & new_n5243;
  assign new_n13914 = ~new_n13909 & ~new_n13913;
  assign new_n13915 = ~new_n13914 & new_n5170;
  assign new_n13916 = ~new_n13905 & ~new_n13915;
  assign new_n13917 = ~new_n13916 & new_n5139;
  assign new_n13918 = ~new_n13895 & ~new_n13917;
  assign new_n13919 = ~new_n5011 & ~new_n13918;
  assign new_n13920 = ~new_n5207 & n3602;
  assign new_n13921 = n3634 & new_n5207;
  assign new_n13922 = ~new_n13920 & ~new_n13921;
  assign new_n13923 = ~new_n5243 & ~new_n13922;
  assign new_n13924 = ~new_n5207 & n3666;
  assign new_n13925 = n3698 & new_n5207;
  assign new_n13926 = ~new_n13924 & ~new_n13925;
  assign new_n13927 = ~new_n13926 & new_n5243;
  assign new_n13928 = ~new_n13923 & ~new_n13927;
  assign new_n13929 = ~new_n5170 & ~new_n13928;
  assign new_n13930 = ~new_n5207 & n3730;
  assign new_n13931 = n3762 & new_n5207;
  assign new_n13932 = ~new_n13930 & ~new_n13931;
  assign new_n13933 = ~new_n5243 & ~new_n13932;
  assign new_n13934 = ~new_n5207 & n3794;
  assign new_n13935 = n3826 & new_n5207;
  assign new_n13936 = ~new_n13934 & ~new_n13935;
  assign new_n13937 = ~new_n13936 & new_n5243;
  assign new_n13938 = ~new_n13933 & ~new_n13937;
  assign new_n13939 = ~new_n13938 & new_n5170;
  assign new_n13940 = ~new_n13929 & ~new_n13939;
  assign new_n13941 = ~new_n5139 & ~new_n13940;
  assign new_n13942 = ~new_n5207 & n3858;
  assign new_n13943 = n3890 & new_n5207;
  assign new_n13944 = ~new_n13942 & ~new_n13943;
  assign new_n13945 = ~new_n5243 & ~new_n13944;
  assign new_n13946 = ~new_n5207 & n3922;
  assign new_n13947 = n3954 & new_n5207;
  assign new_n13948 = ~new_n13946 & ~new_n13947;
  assign new_n13949 = ~new_n13948 & new_n5243;
  assign new_n13950 = ~new_n13945 & ~new_n13949;
  assign new_n13951 = ~new_n5170 & ~new_n13950;
  assign new_n13952 = ~new_n5207 & n3986;
  assign new_n13953 = n4018 & new_n5207;
  assign new_n13954 = ~new_n13952 & ~new_n13953;
  assign new_n13955 = ~new_n5243 & ~new_n13954;
  assign new_n13956 = ~new_n5207 & n4050;
  assign new_n13957 = n4082 & new_n5207;
  assign new_n13958 = ~new_n13956 & ~new_n13957;
  assign new_n13959 = ~new_n13958 & new_n5243;
  assign new_n13960 = ~new_n13955 & ~new_n13959;
  assign new_n13961 = ~new_n13960 & new_n5170;
  assign new_n13962 = ~new_n13951 & ~new_n13961;
  assign new_n13963 = ~new_n13962 & new_n5139;
  assign new_n13964 = ~new_n13941 & ~new_n13963;
  assign new_n13965 = ~new_n13964 & new_n5011;
  assign new_n13966 = ~new_n13919 & ~new_n13965;
  assign new_n13967 = ~new_n13966 & new_n5031;
  assign new_n13968 = ~new_n13873 & ~new_n13967;
  assign new_n13969 = ~new_n5115 & ~new_n13968;
  assign new_n13970 = ~new_n5116 & ~new_n13584;
  assign new_n13971 = ~new_n13969 & ~new_n13970;
  assign new_n13972 = new_n13779 & new_n13971;
  assign new_n13973 = ~new_n9289 & ~new_n13972;
  assign new_n13974 = ~new_n13587 & ~new_n13973;
  assign new_n13975 = ~new_n13972 & new_n8900;
  assign new_n13976 = ~new_n13586 & new_n8901;
  assign new_n13977 = ~new_n13975 & ~new_n13976;
  assign new_n13978 = ~new_n13584 & new_n4150;
  assign new_n13979 = ~new_n5011 & ~new_n9302;
  assign new_n13980 = ~new_n13978 & ~new_n13979;
  assign new_n13981 = new_n13977 & new_n13980;
  assign new_n13982 = new_n13974 & new_n13981;
  assign new_n13983 = ~new_n13982 & new_n8515;
  assign new_n13984 = ~new_n5207 & n2057;
  assign new_n13985 = n2089 & new_n5207;
  assign new_n13986 = ~new_n13984 & ~new_n13985;
  assign new_n13987 = ~new_n5243 & ~new_n13986;
  assign new_n13988 = ~new_n5207 & n2121;
  assign new_n13989 = n2153 & new_n5207;
  assign new_n13990 = ~new_n13988 & ~new_n13989;
  assign new_n13991 = ~new_n13990 & new_n5243;
  assign new_n13992 = ~new_n13987 & ~new_n13991;
  assign new_n13993 = ~new_n5170 & ~new_n13992;
  assign new_n13994 = ~new_n5207 & n2185;
  assign new_n13995 = n2217 & new_n5207;
  assign new_n13996 = ~new_n13994 & ~new_n13995;
  assign new_n13997 = ~new_n5243 & ~new_n13996;
  assign new_n13998 = ~new_n5207 & n2249;
  assign new_n13999 = n2281 & new_n5207;
  assign new_n14000 = ~new_n13998 & ~new_n13999;
  assign new_n14001 = ~new_n14000 & new_n5243;
  assign new_n14002 = ~new_n13997 & ~new_n14001;
  assign new_n14003 = ~new_n14002 & new_n5170;
  assign new_n14004 = ~new_n13993 & ~new_n14003;
  assign new_n14005 = ~new_n5139 & ~new_n14004;
  assign new_n14006 = ~new_n5207 & n2313;
  assign new_n14007 = n2345 & new_n5207;
  assign new_n14008 = ~new_n14006 & ~new_n14007;
  assign new_n14009 = ~new_n5243 & ~new_n14008;
  assign new_n14010 = ~new_n5207 & n2377;
  assign new_n14011 = n2409 & new_n5207;
  assign new_n14012 = ~new_n14010 & ~new_n14011;
  assign new_n14013 = ~new_n14012 & new_n5243;
  assign new_n14014 = ~new_n14009 & ~new_n14013;
  assign new_n14015 = ~new_n5170 & ~new_n14014;
  assign new_n14016 = ~new_n5207 & n2441;
  assign new_n14017 = n2473 & new_n5207;
  assign new_n14018 = ~new_n14016 & ~new_n14017;
  assign new_n14019 = ~new_n5243 & ~new_n14018;
  assign new_n14020 = ~new_n5207 & n2505;
  assign new_n14021 = n2537 & new_n5207;
  assign new_n14022 = ~new_n14020 & ~new_n14021;
  assign new_n14023 = ~new_n14022 & new_n5243;
  assign new_n14024 = ~new_n14019 & ~new_n14023;
  assign new_n14025 = ~new_n14024 & new_n5170;
  assign new_n14026 = ~new_n14015 & ~new_n14025;
  assign new_n14027 = ~new_n14026 & new_n5139;
  assign new_n14028 = ~new_n14005 & ~new_n14027;
  assign new_n14029 = ~new_n5011 & ~new_n14028;
  assign new_n14030 = ~new_n5207 & n2569;
  assign new_n14031 = n2601 & new_n5207;
  assign new_n14032 = ~new_n14030 & ~new_n14031;
  assign new_n14033 = ~new_n5243 & ~new_n14032;
  assign new_n14034 = ~new_n5207 & n2633;
  assign new_n14035 = n2665 & new_n5207;
  assign new_n14036 = ~new_n14034 & ~new_n14035;
  assign new_n14037 = ~new_n14036 & new_n5243;
  assign new_n14038 = ~new_n14033 & ~new_n14037;
  assign new_n14039 = ~new_n5170 & ~new_n14038;
  assign new_n14040 = ~new_n5207 & n2697;
  assign new_n14041 = n2729 & new_n5207;
  assign new_n14042 = ~new_n14040 & ~new_n14041;
  assign new_n14043 = ~new_n5243 & ~new_n14042;
  assign new_n14044 = ~new_n5207 & n2761;
  assign new_n14045 = n2793 & new_n5207;
  assign new_n14046 = ~new_n14044 & ~new_n14045;
  assign new_n14047 = ~new_n14046 & new_n5243;
  assign new_n14048 = ~new_n14043 & ~new_n14047;
  assign new_n14049 = ~new_n14048 & new_n5170;
  assign new_n14050 = ~new_n14039 & ~new_n14049;
  assign new_n14051 = ~new_n5139 & ~new_n14050;
  assign new_n14052 = ~new_n5207 & n2825;
  assign new_n14053 = n2857 & new_n5207;
  assign new_n14054 = ~new_n14052 & ~new_n14053;
  assign new_n14055 = ~new_n5243 & ~new_n14054;
  assign new_n14056 = ~new_n5207 & n2889;
  assign new_n14057 = n2921 & new_n5207;
  assign new_n14058 = ~new_n14056 & ~new_n14057;
  assign new_n14059 = ~new_n14058 & new_n5243;
  assign new_n14060 = ~new_n14055 & ~new_n14059;
  assign new_n14061 = ~new_n5170 & ~new_n14060;
  assign new_n14062 = ~new_n5207 & n2953;
  assign new_n14063 = n2985 & new_n5207;
  assign new_n14064 = ~new_n14062 & ~new_n14063;
  assign new_n14065 = ~new_n5243 & ~new_n14064;
  assign new_n14066 = ~new_n5207 & n3017;
  assign new_n14067 = n3049 & new_n5207;
  assign new_n14068 = ~new_n14066 & ~new_n14067;
  assign new_n14069 = ~new_n14068 & new_n5243;
  assign new_n14070 = ~new_n14065 & ~new_n14069;
  assign new_n14071 = ~new_n14070 & new_n5170;
  assign new_n14072 = ~new_n14061 & ~new_n14071;
  assign new_n14073 = ~new_n14072 & new_n5139;
  assign new_n14074 = ~new_n14051 & ~new_n14073;
  assign new_n14075 = ~new_n14074 & new_n5011;
  assign new_n14076 = ~new_n14029 & ~new_n14075;
  assign new_n14077 = ~new_n5031 & ~new_n14076;
  assign new_n14078 = ~new_n5207 & n3081;
  assign new_n14079 = n3113 & new_n5207;
  assign new_n14080 = ~new_n14078 & ~new_n14079;
  assign new_n14081 = ~new_n5243 & ~new_n14080;
  assign new_n14082 = ~new_n5207 & n3145;
  assign new_n14083 = n3177 & new_n5207;
  assign new_n14084 = ~new_n14082 & ~new_n14083;
  assign new_n14085 = ~new_n14084 & new_n5243;
  assign new_n14086 = ~new_n14081 & ~new_n14085;
  assign new_n14087 = ~new_n5170 & ~new_n14086;
  assign new_n14088 = ~new_n5207 & n3209;
  assign new_n14089 = n3241 & new_n5207;
  assign new_n14090 = ~new_n14088 & ~new_n14089;
  assign new_n14091 = ~new_n5243 & ~new_n14090;
  assign new_n14092 = ~new_n5207 & n3273;
  assign new_n14093 = n3305 & new_n5207;
  assign new_n14094 = ~new_n14092 & ~new_n14093;
  assign new_n14095 = ~new_n14094 & new_n5243;
  assign new_n14096 = ~new_n14091 & ~new_n14095;
  assign new_n14097 = ~new_n14096 & new_n5170;
  assign new_n14098 = ~new_n14087 & ~new_n14097;
  assign new_n14099 = ~new_n5139 & ~new_n14098;
  assign new_n14100 = ~new_n5207 & n3337;
  assign new_n14101 = n3369 & new_n5207;
  assign new_n14102 = ~new_n14100 & ~new_n14101;
  assign new_n14103 = ~new_n5243 & ~new_n14102;
  assign new_n14104 = ~new_n5207 & n3401;
  assign new_n14105 = n3433 & new_n5207;
  assign new_n14106 = ~new_n14104 & ~new_n14105;
  assign new_n14107 = ~new_n14106 & new_n5243;
  assign new_n14108 = ~new_n14103 & ~new_n14107;
  assign new_n14109 = ~new_n5170 & ~new_n14108;
  assign new_n14110 = ~new_n5207 & n3465;
  assign new_n14111 = n3497 & new_n5207;
  assign new_n14112 = ~new_n14110 & ~new_n14111;
  assign new_n14113 = ~new_n5243 & ~new_n14112;
  assign new_n14114 = ~new_n5207 & n3529;
  assign new_n14115 = n3561 & new_n5207;
  assign new_n14116 = ~new_n14114 & ~new_n14115;
  assign new_n14117 = ~new_n14116 & new_n5243;
  assign new_n14118 = ~new_n14113 & ~new_n14117;
  assign new_n14119 = ~new_n14118 & new_n5170;
  assign new_n14120 = ~new_n14109 & ~new_n14119;
  assign new_n14121 = ~new_n14120 & new_n5139;
  assign new_n14122 = ~new_n14099 & ~new_n14121;
  assign new_n14123 = ~new_n5011 & ~new_n14122;
  assign new_n14124 = ~new_n5207 & n3593;
  assign new_n14125 = n3625 & new_n5207;
  assign new_n14126 = ~new_n14124 & ~new_n14125;
  assign new_n14127 = ~new_n5243 & ~new_n14126;
  assign new_n14128 = ~new_n5207 & n3657;
  assign new_n14129 = n3689 & new_n5207;
  assign new_n14130 = ~new_n14128 & ~new_n14129;
  assign new_n14131 = ~new_n14130 & new_n5243;
  assign new_n14132 = ~new_n14127 & ~new_n14131;
  assign new_n14133 = ~new_n5170 & ~new_n14132;
  assign new_n14134 = ~new_n5207 & n3721;
  assign new_n14135 = n3753 & new_n5207;
  assign new_n14136 = ~new_n14134 & ~new_n14135;
  assign new_n14137 = ~new_n5243 & ~new_n14136;
  assign new_n14138 = ~new_n5207 & n3785;
  assign new_n14139 = n3817 & new_n5207;
  assign new_n14140 = ~new_n14138 & ~new_n14139;
  assign new_n14141 = ~new_n14140 & new_n5243;
  assign new_n14142 = ~new_n14137 & ~new_n14141;
  assign new_n14143 = ~new_n14142 & new_n5170;
  assign new_n14144 = ~new_n14133 & ~new_n14143;
  assign new_n14145 = ~new_n5139 & ~new_n14144;
  assign new_n14146 = ~new_n5207 & n3849;
  assign new_n14147 = n3881 & new_n5207;
  assign new_n14148 = ~new_n14146 & ~new_n14147;
  assign new_n14149 = ~new_n5243 & ~new_n14148;
  assign new_n14150 = ~new_n5207 & n3913;
  assign new_n14151 = n3945 & new_n5207;
  assign new_n14152 = ~new_n14150 & ~new_n14151;
  assign new_n14153 = ~new_n14152 & new_n5243;
  assign new_n14154 = ~new_n14149 & ~new_n14153;
  assign new_n14155 = ~new_n5170 & ~new_n14154;
  assign new_n14156 = ~new_n5207 & n3977;
  assign new_n14157 = n4009 & new_n5207;
  assign new_n14158 = ~new_n14156 & ~new_n14157;
  assign new_n14159 = ~new_n5243 & ~new_n14158;
  assign new_n14160 = ~new_n5207 & n4041;
  assign new_n14161 = n4073 & new_n5207;
  assign new_n14162 = ~new_n14160 & ~new_n14161;
  assign new_n14163 = ~new_n14162 & new_n5243;
  assign new_n14164 = ~new_n14159 & ~new_n14163;
  assign new_n14165 = ~new_n14164 & new_n5170;
  assign new_n14166 = ~new_n14155 & ~new_n14165;
  assign new_n14167 = ~new_n14166 & new_n5139;
  assign new_n14168 = ~new_n14145 & ~new_n14167;
  assign new_n14169 = ~new_n14168 & new_n5011;
  assign new_n14170 = ~new_n14123 & ~new_n14169;
  assign new_n14171 = ~new_n14170 & new_n5031;
  assign new_n14172 = ~new_n14077 & ~new_n14171;
  assign new_n14173 = ~new_n5077 & ~new_n14172;
  assign new_n14174 = ~new_n5207 & n2073;
  assign new_n14175 = n2105 & new_n5207;
  assign new_n14176 = ~new_n14174 & ~new_n14175;
  assign new_n14177 = ~new_n5243 & ~new_n14176;
  assign new_n14178 = ~new_n5207 & n2137;
  assign new_n14179 = n2169 & new_n5207;
  assign new_n14180 = ~new_n14178 & ~new_n14179;
  assign new_n14181 = ~new_n14180 & new_n5243;
  assign new_n14182 = ~new_n14177 & ~new_n14181;
  assign new_n14183 = ~new_n5170 & ~new_n14182;
  assign new_n14184 = ~new_n5207 & n2201;
  assign new_n14185 = n2233 & new_n5207;
  assign new_n14186 = ~new_n14184 & ~new_n14185;
  assign new_n14187 = ~new_n5243 & ~new_n14186;
  assign new_n14188 = ~new_n5207 & n2265;
  assign new_n14189 = n2297 & new_n5207;
  assign new_n14190 = ~new_n14188 & ~new_n14189;
  assign new_n14191 = ~new_n14190 & new_n5243;
  assign new_n14192 = ~new_n14187 & ~new_n14191;
  assign new_n14193 = ~new_n14192 & new_n5170;
  assign new_n14194 = ~new_n14183 & ~new_n14193;
  assign new_n14195 = ~new_n5139 & ~new_n14194;
  assign new_n14196 = ~new_n5207 & n2329;
  assign new_n14197 = n2361 & new_n5207;
  assign new_n14198 = ~new_n14196 & ~new_n14197;
  assign new_n14199 = ~new_n5243 & ~new_n14198;
  assign new_n14200 = ~new_n5207 & n2393;
  assign new_n14201 = n2425 & new_n5207;
  assign new_n14202 = ~new_n14200 & ~new_n14201;
  assign new_n14203 = ~new_n14202 & new_n5243;
  assign new_n14204 = ~new_n14199 & ~new_n14203;
  assign new_n14205 = ~new_n5170 & ~new_n14204;
  assign new_n14206 = ~new_n5207 & n2457;
  assign new_n14207 = n2489 & new_n5207;
  assign new_n14208 = ~new_n14206 & ~new_n14207;
  assign new_n14209 = ~new_n5243 & ~new_n14208;
  assign new_n14210 = ~new_n5207 & n2521;
  assign new_n14211 = n2553 & new_n5207;
  assign new_n14212 = ~new_n14210 & ~new_n14211;
  assign new_n14213 = ~new_n14212 & new_n5243;
  assign new_n14214 = ~new_n14209 & ~new_n14213;
  assign new_n14215 = ~new_n14214 & new_n5170;
  assign new_n14216 = ~new_n14205 & ~new_n14215;
  assign new_n14217 = ~new_n14216 & new_n5139;
  assign new_n14218 = ~new_n14195 & ~new_n14217;
  assign new_n14219 = ~new_n5011 & ~new_n14218;
  assign new_n14220 = ~new_n5207 & n2585;
  assign new_n14221 = n2617 & new_n5207;
  assign new_n14222 = ~new_n14220 & ~new_n14221;
  assign new_n14223 = ~new_n5243 & ~new_n14222;
  assign new_n14224 = ~new_n5207 & n2649;
  assign new_n14225 = n2681 & new_n5207;
  assign new_n14226 = ~new_n14224 & ~new_n14225;
  assign new_n14227 = ~new_n14226 & new_n5243;
  assign new_n14228 = ~new_n14223 & ~new_n14227;
  assign new_n14229 = ~new_n5170 & ~new_n14228;
  assign new_n14230 = ~new_n5207 & n2713;
  assign new_n14231 = n2745 & new_n5207;
  assign new_n14232 = ~new_n14230 & ~new_n14231;
  assign new_n14233 = ~new_n5243 & ~new_n14232;
  assign new_n14234 = ~new_n5207 & n2777;
  assign new_n14235 = n2809 & new_n5207;
  assign new_n14236 = ~new_n14234 & ~new_n14235;
  assign new_n14237 = ~new_n14236 & new_n5243;
  assign new_n14238 = ~new_n14233 & ~new_n14237;
  assign new_n14239 = ~new_n14238 & new_n5170;
  assign new_n14240 = ~new_n14229 & ~new_n14239;
  assign new_n14241 = ~new_n5139 & ~new_n14240;
  assign new_n14242 = ~new_n5207 & n2841;
  assign new_n14243 = n2873 & new_n5207;
  assign new_n14244 = ~new_n14242 & ~new_n14243;
  assign new_n14245 = ~new_n5243 & ~new_n14244;
  assign new_n14246 = ~new_n5207 & n2905;
  assign new_n14247 = n2937 & new_n5207;
  assign new_n14248 = ~new_n14246 & ~new_n14247;
  assign new_n14249 = ~new_n14248 & new_n5243;
  assign new_n14250 = ~new_n14245 & ~new_n14249;
  assign new_n14251 = ~new_n5170 & ~new_n14250;
  assign new_n14252 = ~new_n5207 & n2969;
  assign new_n14253 = n3001 & new_n5207;
  assign new_n14254 = ~new_n14252 & ~new_n14253;
  assign new_n14255 = ~new_n5243 & ~new_n14254;
  assign new_n14256 = ~new_n5207 & n3033;
  assign new_n14257 = n3065 & new_n5207;
  assign new_n14258 = ~new_n14256 & ~new_n14257;
  assign new_n14259 = ~new_n14258 & new_n5243;
  assign new_n14260 = ~new_n14255 & ~new_n14259;
  assign new_n14261 = ~new_n14260 & new_n5170;
  assign new_n14262 = ~new_n14251 & ~new_n14261;
  assign new_n14263 = ~new_n14262 & new_n5139;
  assign new_n14264 = ~new_n14241 & ~new_n14263;
  assign new_n14265 = ~new_n14264 & new_n5011;
  assign new_n14266 = ~new_n14219 & ~new_n14265;
  assign new_n14267 = ~new_n5031 & ~new_n14266;
  assign new_n14268 = ~new_n5207 & n3097;
  assign new_n14269 = n3129 & new_n5207;
  assign new_n14270 = ~new_n14268 & ~new_n14269;
  assign new_n14271 = ~new_n5243 & ~new_n14270;
  assign new_n14272 = ~new_n5207 & n3161;
  assign new_n14273 = n3193 & new_n5207;
  assign new_n14274 = ~new_n14272 & ~new_n14273;
  assign new_n14275 = ~new_n14274 & new_n5243;
  assign new_n14276 = ~new_n14271 & ~new_n14275;
  assign new_n14277 = ~new_n5170 & ~new_n14276;
  assign new_n14278 = ~new_n5207 & n3225;
  assign new_n14279 = n3257 & new_n5207;
  assign new_n14280 = ~new_n14278 & ~new_n14279;
  assign new_n14281 = ~new_n5243 & ~new_n14280;
  assign new_n14282 = ~new_n5207 & n3289;
  assign new_n14283 = n3321 & new_n5207;
  assign new_n14284 = ~new_n14282 & ~new_n14283;
  assign new_n14285 = ~new_n14284 & new_n5243;
  assign new_n14286 = ~new_n14281 & ~new_n14285;
  assign new_n14287 = ~new_n14286 & new_n5170;
  assign new_n14288 = ~new_n14277 & ~new_n14287;
  assign new_n14289 = ~new_n5139 & ~new_n14288;
  assign new_n14290 = ~new_n5207 & n3353;
  assign new_n14291 = n3385 & new_n5207;
  assign new_n14292 = ~new_n14290 & ~new_n14291;
  assign new_n14293 = ~new_n5243 & ~new_n14292;
  assign new_n14294 = ~new_n5207 & n3417;
  assign new_n14295 = n3449 & new_n5207;
  assign new_n14296 = ~new_n14294 & ~new_n14295;
  assign new_n14297 = ~new_n14296 & new_n5243;
  assign new_n14298 = ~new_n14293 & ~new_n14297;
  assign new_n14299 = ~new_n5170 & ~new_n14298;
  assign new_n14300 = ~new_n5207 & n3481;
  assign new_n14301 = n3513 & new_n5207;
  assign new_n14302 = ~new_n14300 & ~new_n14301;
  assign new_n14303 = ~new_n5243 & ~new_n14302;
  assign new_n14304 = ~new_n5207 & n3545;
  assign new_n14305 = n3577 & new_n5207;
  assign new_n14306 = ~new_n14304 & ~new_n14305;
  assign new_n14307 = ~new_n14306 & new_n5243;
  assign new_n14308 = ~new_n14303 & ~new_n14307;
  assign new_n14309 = ~new_n14308 & new_n5170;
  assign new_n14310 = ~new_n14299 & ~new_n14309;
  assign new_n14311 = ~new_n14310 & new_n5139;
  assign new_n14312 = ~new_n14289 & ~new_n14311;
  assign new_n14313 = ~new_n5011 & ~new_n14312;
  assign new_n14314 = ~new_n5207 & n3609;
  assign new_n14315 = n3641 & new_n5207;
  assign new_n14316 = ~new_n14314 & ~new_n14315;
  assign new_n14317 = ~new_n5243 & ~new_n14316;
  assign new_n14318 = ~new_n5207 & n3673;
  assign new_n14319 = n3705 & new_n5207;
  assign new_n14320 = ~new_n14318 & ~new_n14319;
  assign new_n14321 = ~new_n14320 & new_n5243;
  assign new_n14322 = ~new_n14317 & ~new_n14321;
  assign new_n14323 = ~new_n5170 & ~new_n14322;
  assign new_n14324 = ~new_n5207 & n3737;
  assign new_n14325 = n3769 & new_n5207;
  assign new_n14326 = ~new_n14324 & ~new_n14325;
  assign new_n14327 = ~new_n5243 & ~new_n14326;
  assign new_n14328 = ~new_n5207 & n3801;
  assign new_n14329 = n3833 & new_n5207;
  assign new_n14330 = ~new_n14328 & ~new_n14329;
  assign new_n14331 = ~new_n14330 & new_n5243;
  assign new_n14332 = ~new_n14327 & ~new_n14331;
  assign new_n14333 = ~new_n14332 & new_n5170;
  assign new_n14334 = ~new_n14323 & ~new_n14333;
  assign new_n14335 = ~new_n5139 & ~new_n14334;
  assign new_n14336 = ~new_n5207 & n3865;
  assign new_n14337 = n3897 & new_n5207;
  assign new_n14338 = ~new_n14336 & ~new_n14337;
  assign new_n14339 = ~new_n5243 & ~new_n14338;
  assign new_n14340 = ~new_n5207 & n3929;
  assign new_n14341 = n3961 & new_n5207;
  assign new_n14342 = ~new_n14340 & ~new_n14341;
  assign new_n14343 = ~new_n14342 & new_n5243;
  assign new_n14344 = ~new_n14339 & ~new_n14343;
  assign new_n14345 = ~new_n5170 & ~new_n14344;
  assign new_n14346 = ~new_n5207 & n3993;
  assign new_n14347 = n4025 & new_n5207;
  assign new_n14348 = ~new_n14346 & ~new_n14347;
  assign new_n14349 = ~new_n5243 & ~new_n14348;
  assign new_n14350 = ~new_n5207 & n4057;
  assign new_n14351 = n4089 & new_n5207;
  assign new_n14352 = ~new_n14350 & ~new_n14351;
  assign new_n14353 = ~new_n14352 & new_n5243;
  assign new_n14354 = ~new_n14349 & ~new_n14353;
  assign new_n14355 = ~new_n14354 & new_n5170;
  assign new_n14356 = ~new_n14345 & ~new_n14355;
  assign new_n14357 = ~new_n14356 & new_n5139;
  assign new_n14358 = ~new_n14335 & ~new_n14357;
  assign new_n14359 = ~new_n14358 & new_n5011;
  assign new_n14360 = ~new_n14313 & ~new_n14359;
  assign new_n14361 = ~new_n14360 & new_n5031;
  assign new_n14362 = ~new_n14267 & ~new_n14361;
  assign new_n14363 = ~new_n14362 & new_n5077;
  assign new_n14364 = ~new_n14173 & ~new_n14363;
  assign new_n14365 = ~new_n14364 & new_n8902;
  assign new_n14366 = ~new_n5207 & n2049;
  assign new_n14367 = n2081 & new_n5207;
  assign new_n14368 = ~new_n14366 & ~new_n14367;
  assign new_n14369 = ~new_n5243 & ~new_n14368;
  assign new_n14370 = ~new_n5207 & n2113;
  assign new_n14371 = n2145 & new_n5207;
  assign new_n14372 = ~new_n14370 & ~new_n14371;
  assign new_n14373 = ~new_n14372 & new_n5243;
  assign new_n14374 = ~new_n14369 & ~new_n14373;
  assign new_n14375 = ~new_n5170 & ~new_n14374;
  assign new_n14376 = ~new_n5207 & n2177;
  assign new_n14377 = n2209 & new_n5207;
  assign new_n14378 = ~new_n14376 & ~new_n14377;
  assign new_n14379 = ~new_n5243 & ~new_n14378;
  assign new_n14380 = ~new_n5207 & n2241;
  assign new_n14381 = n2273 & new_n5207;
  assign new_n14382 = ~new_n14380 & ~new_n14381;
  assign new_n14383 = ~new_n14382 & new_n5243;
  assign new_n14384 = ~new_n14379 & ~new_n14383;
  assign new_n14385 = ~new_n14384 & new_n5170;
  assign new_n14386 = ~new_n14375 & ~new_n14385;
  assign new_n14387 = ~new_n5139 & ~new_n14386;
  assign new_n14388 = ~new_n5207 & n2305;
  assign new_n14389 = n2337 & new_n5207;
  assign new_n14390 = ~new_n14388 & ~new_n14389;
  assign new_n14391 = ~new_n5243 & ~new_n14390;
  assign new_n14392 = ~new_n5207 & n2369;
  assign new_n14393 = n2401 & new_n5207;
  assign new_n14394 = ~new_n14392 & ~new_n14393;
  assign new_n14395 = ~new_n14394 & new_n5243;
  assign new_n14396 = ~new_n14391 & ~new_n14395;
  assign new_n14397 = ~new_n5170 & ~new_n14396;
  assign new_n14398 = ~new_n5207 & n2433;
  assign new_n14399 = n2465 & new_n5207;
  assign new_n14400 = ~new_n14398 & ~new_n14399;
  assign new_n14401 = ~new_n5243 & ~new_n14400;
  assign new_n14402 = ~new_n5207 & n2497;
  assign new_n14403 = n2529 & new_n5207;
  assign new_n14404 = ~new_n14402 & ~new_n14403;
  assign new_n14405 = ~new_n14404 & new_n5243;
  assign new_n14406 = ~new_n14401 & ~new_n14405;
  assign new_n14407 = ~new_n14406 & new_n5170;
  assign new_n14408 = ~new_n14397 & ~new_n14407;
  assign new_n14409 = ~new_n14408 & new_n5139;
  assign new_n14410 = ~new_n14387 & ~new_n14409;
  assign new_n14411 = ~new_n5011 & ~new_n14410;
  assign new_n14412 = ~new_n5207 & n2561;
  assign new_n14413 = n2593 & new_n5207;
  assign new_n14414 = ~new_n14412 & ~new_n14413;
  assign new_n14415 = ~new_n5243 & ~new_n14414;
  assign new_n14416 = ~new_n5207 & n2625;
  assign new_n14417 = n2657 & new_n5207;
  assign new_n14418 = ~new_n14416 & ~new_n14417;
  assign new_n14419 = ~new_n14418 & new_n5243;
  assign new_n14420 = ~new_n14415 & ~new_n14419;
  assign new_n14421 = ~new_n5170 & ~new_n14420;
  assign new_n14422 = ~new_n5207 & n2689;
  assign new_n14423 = n2721 & new_n5207;
  assign new_n14424 = ~new_n14422 & ~new_n14423;
  assign new_n14425 = ~new_n5243 & ~new_n14424;
  assign new_n14426 = ~new_n5207 & n2753;
  assign new_n14427 = n2785 & new_n5207;
  assign new_n14428 = ~new_n14426 & ~new_n14427;
  assign new_n14429 = ~new_n14428 & new_n5243;
  assign new_n14430 = ~new_n14425 & ~new_n14429;
  assign new_n14431 = ~new_n14430 & new_n5170;
  assign new_n14432 = ~new_n14421 & ~new_n14431;
  assign new_n14433 = ~new_n5139 & ~new_n14432;
  assign new_n14434 = ~new_n5207 & n2817;
  assign new_n14435 = n2849 & new_n5207;
  assign new_n14436 = ~new_n14434 & ~new_n14435;
  assign new_n14437 = ~new_n5243 & ~new_n14436;
  assign new_n14438 = ~new_n5207 & n2881;
  assign new_n14439 = n2913 & new_n5207;
  assign new_n14440 = ~new_n14438 & ~new_n14439;
  assign new_n14441 = ~new_n14440 & new_n5243;
  assign new_n14442 = ~new_n14437 & ~new_n14441;
  assign new_n14443 = ~new_n5170 & ~new_n14442;
  assign new_n14444 = ~new_n5207 & n2945;
  assign new_n14445 = n2977 & new_n5207;
  assign new_n14446 = ~new_n14444 & ~new_n14445;
  assign new_n14447 = ~new_n5243 & ~new_n14446;
  assign new_n14448 = ~new_n5207 & n3009;
  assign new_n14449 = n3041 & new_n5207;
  assign new_n14450 = ~new_n14448 & ~new_n14449;
  assign new_n14451 = ~new_n14450 & new_n5243;
  assign new_n14452 = ~new_n14447 & ~new_n14451;
  assign new_n14453 = ~new_n14452 & new_n5170;
  assign new_n14454 = ~new_n14443 & ~new_n14453;
  assign new_n14455 = ~new_n14454 & new_n5139;
  assign new_n14456 = ~new_n14433 & ~new_n14455;
  assign new_n14457 = ~new_n14456 & new_n5011;
  assign new_n14458 = ~new_n14411 & ~new_n14457;
  assign new_n14459 = ~new_n5031 & ~new_n14458;
  assign new_n14460 = ~new_n5207 & n3073;
  assign new_n14461 = n3105 & new_n5207;
  assign new_n14462 = ~new_n14460 & ~new_n14461;
  assign new_n14463 = ~new_n5243 & ~new_n14462;
  assign new_n14464 = ~new_n5207 & n3137;
  assign new_n14465 = n3169 & new_n5207;
  assign new_n14466 = ~new_n14464 & ~new_n14465;
  assign new_n14467 = ~new_n14466 & new_n5243;
  assign new_n14468 = ~new_n14463 & ~new_n14467;
  assign new_n14469 = ~new_n5170 & ~new_n14468;
  assign new_n14470 = ~new_n5207 & n3201;
  assign new_n14471 = n3233 & new_n5207;
  assign new_n14472 = ~new_n14470 & ~new_n14471;
  assign new_n14473 = ~new_n5243 & ~new_n14472;
  assign new_n14474 = ~new_n5207 & n3265;
  assign new_n14475 = n3297 & new_n5207;
  assign new_n14476 = ~new_n14474 & ~new_n14475;
  assign new_n14477 = ~new_n14476 & new_n5243;
  assign new_n14478 = ~new_n14473 & ~new_n14477;
  assign new_n14479 = ~new_n14478 & new_n5170;
  assign new_n14480 = ~new_n14469 & ~new_n14479;
  assign new_n14481 = ~new_n5139 & ~new_n14480;
  assign new_n14482 = ~new_n5207 & n3329;
  assign new_n14483 = n3361 & new_n5207;
  assign new_n14484 = ~new_n14482 & ~new_n14483;
  assign new_n14485 = ~new_n5243 & ~new_n14484;
  assign new_n14486 = ~new_n5207 & n3393;
  assign new_n14487 = n3425 & new_n5207;
  assign new_n14488 = ~new_n14486 & ~new_n14487;
  assign new_n14489 = ~new_n14488 & new_n5243;
  assign new_n14490 = ~new_n14485 & ~new_n14489;
  assign new_n14491 = ~new_n5170 & ~new_n14490;
  assign new_n14492 = ~new_n5207 & n3457;
  assign new_n14493 = n3489 & new_n5207;
  assign new_n14494 = ~new_n14492 & ~new_n14493;
  assign new_n14495 = ~new_n5243 & ~new_n14494;
  assign new_n14496 = ~new_n5207 & n3521;
  assign new_n14497 = n3553 & new_n5207;
  assign new_n14498 = ~new_n14496 & ~new_n14497;
  assign new_n14499 = ~new_n14498 & new_n5243;
  assign new_n14500 = ~new_n14495 & ~new_n14499;
  assign new_n14501 = ~new_n14500 & new_n5170;
  assign new_n14502 = ~new_n14491 & ~new_n14501;
  assign new_n14503 = ~new_n14502 & new_n5139;
  assign new_n14504 = ~new_n14481 & ~new_n14503;
  assign new_n14505 = ~new_n5011 & ~new_n14504;
  assign new_n14506 = ~new_n5207 & n3585;
  assign new_n14507 = n3617 & new_n5207;
  assign new_n14508 = ~new_n14506 & ~new_n14507;
  assign new_n14509 = ~new_n5243 & ~new_n14508;
  assign new_n14510 = ~new_n5207 & n3649;
  assign new_n14511 = n3681 & new_n5207;
  assign new_n14512 = ~new_n14510 & ~new_n14511;
  assign new_n14513 = ~new_n14512 & new_n5243;
  assign new_n14514 = ~new_n14509 & ~new_n14513;
  assign new_n14515 = ~new_n5170 & ~new_n14514;
  assign new_n14516 = ~new_n5207 & n3713;
  assign new_n14517 = n3745 & new_n5207;
  assign new_n14518 = ~new_n14516 & ~new_n14517;
  assign new_n14519 = ~new_n5243 & ~new_n14518;
  assign new_n14520 = ~new_n5207 & n3777;
  assign new_n14521 = n3809 & new_n5207;
  assign new_n14522 = ~new_n14520 & ~new_n14521;
  assign new_n14523 = ~new_n14522 & new_n5243;
  assign new_n14524 = ~new_n14519 & ~new_n14523;
  assign new_n14525 = ~new_n14524 & new_n5170;
  assign new_n14526 = ~new_n14515 & ~new_n14525;
  assign new_n14527 = ~new_n5139 & ~new_n14526;
  assign new_n14528 = ~new_n5207 & n3841;
  assign new_n14529 = n3873 & new_n5207;
  assign new_n14530 = ~new_n14528 & ~new_n14529;
  assign new_n14531 = ~new_n5243 & ~new_n14530;
  assign new_n14532 = ~new_n5207 & n3905;
  assign new_n14533 = n3937 & new_n5207;
  assign new_n14534 = ~new_n14532 & ~new_n14533;
  assign new_n14535 = ~new_n14534 & new_n5243;
  assign new_n14536 = ~new_n14531 & ~new_n14535;
  assign new_n14537 = ~new_n5170 & ~new_n14536;
  assign new_n14538 = ~new_n5207 & n3969;
  assign new_n14539 = n4001 & new_n5207;
  assign new_n14540 = ~new_n14538 & ~new_n14539;
  assign new_n14541 = ~new_n5243 & ~new_n14540;
  assign new_n14542 = ~new_n5207 & n4033;
  assign new_n14543 = n4065 & new_n5207;
  assign new_n14544 = ~new_n14542 & ~new_n14543;
  assign new_n14545 = ~new_n14544 & new_n5243;
  assign new_n14546 = ~new_n14541 & ~new_n14545;
  assign new_n14547 = ~new_n14546 & new_n5170;
  assign new_n14548 = ~new_n14537 & ~new_n14547;
  assign new_n14549 = ~new_n14548 & new_n5139;
  assign new_n14550 = ~new_n14527 & ~new_n14549;
  assign new_n14551 = ~new_n14550 & new_n5011;
  assign new_n14552 = ~new_n14505 & ~new_n14551;
  assign new_n14553 = ~new_n14552 & new_n5031;
  assign new_n14554 = ~new_n14459 & ~new_n14553;
  assign new_n14555 = ~new_n14554 & new_n5114;
  assign new_n14556 = ~new_n5462 & ~new_n14172;
  assign new_n14557 = ~new_n14555 & ~new_n14556;
  assign new_n14558 = ~new_n5207 & n2065;
  assign new_n14559 = n2097 & new_n5207;
  assign new_n14560 = ~new_n14558 & ~new_n14559;
  assign new_n14561 = ~new_n5243 & ~new_n14560;
  assign new_n14562 = ~new_n5207 & n2129;
  assign new_n14563 = n2161 & new_n5207;
  assign new_n14564 = ~new_n14562 & ~new_n14563;
  assign new_n14565 = ~new_n14564 & new_n5243;
  assign new_n14566 = ~new_n14561 & ~new_n14565;
  assign new_n14567 = ~new_n5170 & ~new_n14566;
  assign new_n14568 = ~new_n5207 & n2193;
  assign new_n14569 = n2225 & new_n5207;
  assign new_n14570 = ~new_n14568 & ~new_n14569;
  assign new_n14571 = ~new_n5243 & ~new_n14570;
  assign new_n14572 = ~new_n5207 & n2257;
  assign new_n14573 = n2289 & new_n5207;
  assign new_n14574 = ~new_n14572 & ~new_n14573;
  assign new_n14575 = ~new_n14574 & new_n5243;
  assign new_n14576 = ~new_n14571 & ~new_n14575;
  assign new_n14577 = ~new_n14576 & new_n5170;
  assign new_n14578 = ~new_n14567 & ~new_n14577;
  assign new_n14579 = ~new_n5139 & ~new_n14578;
  assign new_n14580 = ~new_n5207 & n2321;
  assign new_n14581 = n2353 & new_n5207;
  assign new_n14582 = ~new_n14580 & ~new_n14581;
  assign new_n14583 = ~new_n5243 & ~new_n14582;
  assign new_n14584 = ~new_n5207 & n2385;
  assign new_n14585 = n2417 & new_n5207;
  assign new_n14586 = ~new_n14584 & ~new_n14585;
  assign new_n14587 = ~new_n14586 & new_n5243;
  assign new_n14588 = ~new_n14583 & ~new_n14587;
  assign new_n14589 = ~new_n5170 & ~new_n14588;
  assign new_n14590 = ~new_n5207 & n2449;
  assign new_n14591 = n2481 & new_n5207;
  assign new_n14592 = ~new_n14590 & ~new_n14591;
  assign new_n14593 = ~new_n5243 & ~new_n14592;
  assign new_n14594 = ~new_n5207 & n2513;
  assign new_n14595 = n2545 & new_n5207;
  assign new_n14596 = ~new_n14594 & ~new_n14595;
  assign new_n14597 = ~new_n14596 & new_n5243;
  assign new_n14598 = ~new_n14593 & ~new_n14597;
  assign new_n14599 = ~new_n14598 & new_n5170;
  assign new_n14600 = ~new_n14589 & ~new_n14599;
  assign new_n14601 = ~new_n14600 & new_n5139;
  assign new_n14602 = ~new_n14579 & ~new_n14601;
  assign new_n14603 = ~new_n5011 & ~new_n14602;
  assign new_n14604 = ~new_n5207 & n2577;
  assign new_n14605 = n2609 & new_n5207;
  assign new_n14606 = ~new_n14604 & ~new_n14605;
  assign new_n14607 = ~new_n5243 & ~new_n14606;
  assign new_n14608 = ~new_n5207 & n2641;
  assign new_n14609 = n2673 & new_n5207;
  assign new_n14610 = ~new_n14608 & ~new_n14609;
  assign new_n14611 = ~new_n14610 & new_n5243;
  assign new_n14612 = ~new_n14607 & ~new_n14611;
  assign new_n14613 = ~new_n5170 & ~new_n14612;
  assign new_n14614 = ~new_n5207 & n2705;
  assign new_n14615 = n2737 & new_n5207;
  assign new_n14616 = ~new_n14614 & ~new_n14615;
  assign new_n14617 = ~new_n5243 & ~new_n14616;
  assign new_n14618 = ~new_n5207 & n2769;
  assign new_n14619 = n2801 & new_n5207;
  assign new_n14620 = ~new_n14618 & ~new_n14619;
  assign new_n14621 = ~new_n14620 & new_n5243;
  assign new_n14622 = ~new_n14617 & ~new_n14621;
  assign new_n14623 = ~new_n14622 & new_n5170;
  assign new_n14624 = ~new_n14613 & ~new_n14623;
  assign new_n14625 = ~new_n5139 & ~new_n14624;
  assign new_n14626 = ~new_n5207 & n2833;
  assign new_n14627 = n2865 & new_n5207;
  assign new_n14628 = ~new_n14626 & ~new_n14627;
  assign new_n14629 = ~new_n5243 & ~new_n14628;
  assign new_n14630 = ~new_n5207 & n2897;
  assign new_n14631 = n2929 & new_n5207;
  assign new_n14632 = ~new_n14630 & ~new_n14631;
  assign new_n14633 = ~new_n14632 & new_n5243;
  assign new_n14634 = ~new_n14629 & ~new_n14633;
  assign new_n14635 = ~new_n5170 & ~new_n14634;
  assign new_n14636 = ~new_n5207 & n2961;
  assign new_n14637 = n2993 & new_n5207;
  assign new_n14638 = ~new_n14636 & ~new_n14637;
  assign new_n14639 = ~new_n5243 & ~new_n14638;
  assign new_n14640 = ~new_n5207 & n3025;
  assign new_n14641 = n3057 & new_n5207;
  assign new_n14642 = ~new_n14640 & ~new_n14641;
  assign new_n14643 = ~new_n14642 & new_n5243;
  assign new_n14644 = ~new_n14639 & ~new_n14643;
  assign new_n14645 = ~new_n14644 & new_n5170;
  assign new_n14646 = ~new_n14635 & ~new_n14645;
  assign new_n14647 = ~new_n14646 & new_n5139;
  assign new_n14648 = ~new_n14625 & ~new_n14647;
  assign new_n14649 = ~new_n14648 & new_n5011;
  assign new_n14650 = ~new_n14603 & ~new_n14649;
  assign new_n14651 = ~new_n5031 & ~new_n14650;
  assign new_n14652 = ~new_n5207 & n3089;
  assign new_n14653 = n3121 & new_n5207;
  assign new_n14654 = ~new_n14652 & ~new_n14653;
  assign new_n14655 = ~new_n5243 & ~new_n14654;
  assign new_n14656 = ~new_n5207 & n3153;
  assign new_n14657 = n3185 & new_n5207;
  assign new_n14658 = ~new_n14656 & ~new_n14657;
  assign new_n14659 = ~new_n14658 & new_n5243;
  assign new_n14660 = ~new_n14655 & ~new_n14659;
  assign new_n14661 = ~new_n5170 & ~new_n14660;
  assign new_n14662 = ~new_n5207 & n3217;
  assign new_n14663 = n3249 & new_n5207;
  assign new_n14664 = ~new_n14662 & ~new_n14663;
  assign new_n14665 = ~new_n5243 & ~new_n14664;
  assign new_n14666 = ~new_n5207 & n3281;
  assign new_n14667 = n3313 & new_n5207;
  assign new_n14668 = ~new_n14666 & ~new_n14667;
  assign new_n14669 = ~new_n14668 & new_n5243;
  assign new_n14670 = ~new_n14665 & ~new_n14669;
  assign new_n14671 = ~new_n14670 & new_n5170;
  assign new_n14672 = ~new_n14661 & ~new_n14671;
  assign new_n14673 = ~new_n5139 & ~new_n14672;
  assign new_n14674 = ~new_n5207 & n3345;
  assign new_n14675 = n3377 & new_n5207;
  assign new_n14676 = ~new_n14674 & ~new_n14675;
  assign new_n14677 = ~new_n5243 & ~new_n14676;
  assign new_n14678 = ~new_n5207 & n3409;
  assign new_n14679 = n3441 & new_n5207;
  assign new_n14680 = ~new_n14678 & ~new_n14679;
  assign new_n14681 = ~new_n14680 & new_n5243;
  assign new_n14682 = ~new_n14677 & ~new_n14681;
  assign new_n14683 = ~new_n5170 & ~new_n14682;
  assign new_n14684 = ~new_n5207 & n3473;
  assign new_n14685 = n3505 & new_n5207;
  assign new_n14686 = ~new_n14684 & ~new_n14685;
  assign new_n14687 = ~new_n5243 & ~new_n14686;
  assign new_n14688 = ~new_n5207 & n3537;
  assign new_n14689 = n3569 & new_n5207;
  assign new_n14690 = ~new_n14688 & ~new_n14689;
  assign new_n14691 = ~new_n14690 & new_n5243;
  assign new_n14692 = ~new_n14687 & ~new_n14691;
  assign new_n14693 = ~new_n14692 & new_n5170;
  assign new_n14694 = ~new_n14683 & ~new_n14693;
  assign new_n14695 = ~new_n14694 & new_n5139;
  assign new_n14696 = ~new_n14673 & ~new_n14695;
  assign new_n14697 = ~new_n5011 & ~new_n14696;
  assign new_n14698 = ~new_n5207 & n3601;
  assign new_n14699 = n3633 & new_n5207;
  assign new_n14700 = ~new_n14698 & ~new_n14699;
  assign new_n14701 = ~new_n5243 & ~new_n14700;
  assign new_n14702 = ~new_n5207 & n3665;
  assign new_n14703 = n3697 & new_n5207;
  assign new_n14704 = ~new_n14702 & ~new_n14703;
  assign new_n14705 = ~new_n14704 & new_n5243;
  assign new_n14706 = ~new_n14701 & ~new_n14705;
  assign new_n14707 = ~new_n5170 & ~new_n14706;
  assign new_n14708 = ~new_n5207 & n3729;
  assign new_n14709 = n3761 & new_n5207;
  assign new_n14710 = ~new_n14708 & ~new_n14709;
  assign new_n14711 = ~new_n5243 & ~new_n14710;
  assign new_n14712 = ~new_n5207 & n3793;
  assign new_n14713 = n3825 & new_n5207;
  assign new_n14714 = ~new_n14712 & ~new_n14713;
  assign new_n14715 = ~new_n14714 & new_n5243;
  assign new_n14716 = ~new_n14711 & ~new_n14715;
  assign new_n14717 = ~new_n14716 & new_n5170;
  assign new_n14718 = ~new_n14707 & ~new_n14717;
  assign new_n14719 = ~new_n5139 & ~new_n14718;
  assign new_n14720 = ~new_n5207 & n3857;
  assign new_n14721 = n3889 & new_n5207;
  assign new_n14722 = ~new_n14720 & ~new_n14721;
  assign new_n14723 = ~new_n5243 & ~new_n14722;
  assign new_n14724 = ~new_n5207 & n3921;
  assign new_n14725 = n3953 & new_n5207;
  assign new_n14726 = ~new_n14724 & ~new_n14725;
  assign new_n14727 = ~new_n14726 & new_n5243;
  assign new_n14728 = ~new_n14723 & ~new_n14727;
  assign new_n14729 = ~new_n5170 & ~new_n14728;
  assign new_n14730 = ~new_n5207 & n3985;
  assign new_n14731 = n4017 & new_n5207;
  assign new_n14732 = ~new_n14730 & ~new_n14731;
  assign new_n14733 = ~new_n5243 & ~new_n14732;
  assign new_n14734 = ~new_n5207 & n4049;
  assign new_n14735 = n4081 & new_n5207;
  assign new_n14736 = ~new_n14734 & ~new_n14735;
  assign new_n14737 = ~new_n14736 & new_n5243;
  assign new_n14738 = ~new_n14733 & ~new_n14737;
  assign new_n14739 = ~new_n14738 & new_n5170;
  assign new_n14740 = ~new_n14729 & ~new_n14739;
  assign new_n14741 = ~new_n14740 & new_n5139;
  assign new_n14742 = ~new_n14719 & ~new_n14741;
  assign new_n14743 = ~new_n14742 & new_n5011;
  assign new_n14744 = ~new_n14697 & ~new_n14743;
  assign new_n14745 = ~new_n14744 & new_n5031;
  assign new_n14746 = ~new_n14651 & ~new_n14745;
  assign new_n14747 = ~new_n5115 & ~new_n14746;
  assign new_n14748 = ~new_n5116 & ~new_n14362;
  assign new_n14749 = ~new_n14747 & ~new_n14748;
  assign new_n14750 = new_n14557 & new_n14749;
  assign new_n14751 = ~new_n9289 & ~new_n14750;
  assign new_n14752 = ~new_n14365 & ~new_n14751;
  assign new_n14753 = ~new_n14750 & new_n8900;
  assign new_n14754 = ~new_n14364 & new_n8901;
  assign new_n14755 = ~new_n14753 & ~new_n14754;
  assign new_n14756 = ~new_n14362 & new_n4150;
  assign new_n14757 = ~new_n5031 & ~new_n9302;
  assign new_n14758 = ~new_n14756 & ~new_n14757;
  assign new_n14759 = new_n14755 & new_n14758;
  assign new_n14760 = new_n14752 & new_n14759;
  assign new_n14761 = ~new_n14760 & new_n8515;
  assign new_n14762 = ~new_n4964 & ~new_n9302;
  assign new_n14763 = ~new_n14362 & new_n8900;
  assign new_n14764 = ~new_n14762 & ~new_n14763;
  assign new_n14765 = ~new_n9284 & new_n4150;
  assign new_n14766 = ~new_n14765 & new_n14764;
  assign new_n14767 = ~new_n5077 & ~new_n9092;
  assign new_n14768 = ~new_n9284 & new_n5077;
  assign new_n14769 = ~new_n14767 & ~new_n14768;
  assign new_n14770 = ~new_n14769 & new_n8898;
  assign new_n14771 = ~new_n14770 & new_n14766;
  assign new_n14772 = ~new_n14771 & new_n8515;
  assign new_n14773 = ~new_n4988 & ~new_n9302;
  assign new_n14774 = ~new_n14763 & ~new_n14773;
  assign new_n14775 = ~new_n10074 & new_n4150;
  assign new_n14776 = ~new_n14775 & new_n14774;
  assign new_n14777 = ~new_n5077 & ~new_n9882;
  assign new_n14778 = ~new_n10074 & new_n5077;
  assign new_n14779 = ~new_n14777 & ~new_n14778;
  assign new_n14780 = ~new_n14779 & new_n8898;
  assign new_n14781 = ~new_n14780 & new_n14776;
  assign new_n14782 = ~new_n14781 & new_n8515;
  assign new_n14783 = ~new_n4915 & ~new_n9302;
  assign new_n14784 = ~new_n14763 & ~new_n14783;
  assign new_n14785 = ~new_n10855 & new_n4150;
  assign new_n14786 = ~new_n14785 & new_n14784;
  assign new_n14787 = ~new_n5077 & ~new_n10663;
  assign new_n14788 = ~new_n10855 & new_n5077;
  assign new_n14789 = ~new_n14787 & ~new_n14788;
  assign new_n14790 = ~new_n14789 & new_n8898;
  assign new_n14791 = ~new_n14790 & new_n14786;
  assign new_n14792 = ~new_n14791 & new_n8515;
  assign new_n14793 = ~new_n4939 & ~new_n9302;
  assign new_n14794 = ~new_n14763 & ~new_n14793;
  assign new_n14795 = ~new_n11634 & new_n4150;
  assign new_n14796 = ~new_n14795 & new_n14794;
  assign new_n14797 = ~new_n5077 & ~new_n11442;
  assign new_n14798 = ~new_n11634 & new_n5077;
  assign new_n14799 = ~new_n14797 & ~new_n14798;
  assign new_n14800 = ~new_n14799 & new_n8898;
  assign new_n14801 = ~new_n14800 & new_n14796;
  assign new_n14802 = ~new_n14801 & new_n8515;
  assign new_n14803 = ~new_n4866 & ~new_n9302;
  assign new_n14804 = ~new_n14763 & ~new_n14803;
  assign new_n14805 = ~new_n12412 & new_n4150;
  assign new_n14806 = ~new_n14805 & new_n14804;
  assign new_n14807 = ~new_n5077 & ~new_n12220;
  assign new_n14808 = ~new_n12412 & new_n5077;
  assign new_n14809 = ~new_n14807 & ~new_n14808;
  assign new_n14810 = ~new_n14809 & new_n8898;
  assign new_n14811 = ~new_n14810 & new_n14806;
  assign new_n14812 = ~new_n14811 & new_n8515;
  assign new_n14813 = ~new_n4889 & ~new_n9302;
  assign new_n14814 = ~new_n14763 & ~new_n14813;
  assign new_n14815 = ~new_n13190 & new_n4150;
  assign new_n14816 = ~new_n14815 & new_n14814;
  assign new_n14817 = ~new_n5077 & ~new_n12998;
  assign new_n14818 = ~new_n13190 & new_n5077;
  assign new_n14819 = ~new_n14817 & ~new_n14818;
  assign new_n14820 = ~new_n14819 & new_n8898;
  assign new_n14821 = ~new_n14820 & new_n14816;
  assign new_n14822 = ~new_n14821 & new_n8515;
  assign new_n14823 = ~new_n4818 & ~new_n9302;
  assign new_n14824 = ~new_n14763 & ~new_n14823;
  assign new_n14825 = ~new_n13968 & new_n4150;
  assign new_n14826 = ~new_n14825 & new_n14824;
  assign new_n14827 = ~new_n5077 & ~new_n13776;
  assign new_n14828 = ~new_n13968 & new_n5077;
  assign new_n14829 = ~new_n14827 & ~new_n14828;
  assign new_n14830 = ~new_n14829 & new_n8898;
  assign new_n14831 = ~new_n14830 & new_n14826;
  assign new_n14832 = ~new_n14831 & new_n8515;
  assign new_n14833 = ~new_n4842 & ~new_n9302;
  assign new_n14834 = ~new_n14763 & ~new_n14833;
  assign new_n14835 = ~new_n14746 & new_n4150;
  assign new_n14836 = ~new_n14835 & new_n14834;
  assign new_n14837 = ~new_n5077 & ~new_n14554;
  assign new_n14838 = ~new_n14746 & new_n5077;
  assign new_n14839 = ~new_n14837 & ~new_n14838;
  assign new_n14840 = ~new_n14839 & new_n8898;
  assign new_n14841 = ~new_n14840 & new_n14836;
  assign new_n14842 = ~new_n14841 & new_n8515;
  assign new_n14843 = new_n14838 ^ new_n8895;
  assign new_n14844 = new_n8901 & new_n14843;
  assign new_n14845 = ~new_n14763 & ~new_n14844;
  assign new_n14846 = n2048 & new_n4138;
  assign new_n14847 = ~new_n14846 & new_n14845;
  assign new_n14848 = ~new_n4772 & ~new_n9302;
  assign new_n14849 = ~new_n8894 & new_n4150;
  assign new_n14850 = ~new_n14848 & ~new_n14849;
  assign new_n14851 = new_n14847 & new_n14850;
  assign new_n14852 = ~new_n14851 & new_n8515;
  assign new_n14853 = n2047 & new_n4138;
  assign new_n14854 = ~new_n14853 & new_n14845;
  assign new_n14855 = ~new_n4785 & ~new_n9302;
  assign new_n14856 = ~new_n9500 & new_n4150;
  assign new_n14857 = ~new_n14855 & ~new_n14856;
  assign new_n14858 = new_n14854 & new_n14857;
  assign new_n14859 = ~new_n14858 & new_n8515;
  assign new_n14860 = n2046 & new_n4138;
  assign new_n14861 = ~new_n14860 & new_n14845;
  assign new_n14862 = ~new_n4747 & ~new_n9302;
  assign new_n14863 = ~new_n10281 & new_n4150;
  assign new_n14864 = ~new_n14862 & ~new_n14863;
  assign new_n14865 = new_n14861 & new_n14864;
  assign new_n14866 = ~new_n14865 & new_n8515;
  assign new_n14867 = n2045 & new_n4138;
  assign new_n14868 = ~new_n14867 & new_n14845;
  assign new_n14869 = ~new_n4759 & ~new_n9302;
  assign new_n14870 = ~new_n11060 & new_n4150;
  assign new_n14871 = ~new_n14869 & ~new_n14870;
  assign new_n14872 = new_n14868 & new_n14871;
  assign new_n14873 = ~new_n14872 & new_n8515;
  assign new_n14874 = n2044 & new_n4138;
  assign new_n14875 = ~new_n14874 & new_n14845;
  assign new_n14876 = ~new_n4717 & ~new_n9302;
  assign new_n14877 = ~new_n11838 & new_n4150;
  assign new_n14878 = ~new_n14876 & ~new_n14877;
  assign new_n14879 = new_n14875 & new_n14878;
  assign new_n14880 = ~new_n14879 & new_n8515;
  assign new_n14881 = n2043 & new_n4138;
  assign new_n14882 = ~new_n14881 & new_n14845;
  assign new_n14883 = ~new_n4731 & ~new_n9302;
  assign new_n14884 = ~new_n12616 & new_n4150;
  assign new_n14885 = ~new_n14883 & ~new_n14884;
  assign new_n14886 = new_n14882 & new_n14885;
  assign new_n14887 = ~new_n14886 & new_n8515;
  assign new_n14888 = n2042 & new_n4138;
  assign new_n14889 = ~new_n14888 & new_n14845;
  assign new_n14890 = ~new_n4685 & ~new_n9302;
  assign new_n14891 = ~new_n13394 & new_n4150;
  assign new_n14892 = ~new_n14890 & ~new_n14891;
  assign new_n14893 = new_n14889 & new_n14892;
  assign new_n14894 = ~new_n14893 & new_n8515;
  assign new_n14895 = n2041 & new_n4138;
  assign new_n14896 = ~new_n14895 & new_n14845;
  assign new_n14897 = ~new_n4699 & ~new_n9302;
  assign new_n14898 = ~new_n14172 & new_n4150;
  assign new_n14899 = ~new_n14897 & ~new_n14898;
  assign new_n14900 = new_n14896 & new_n14899;
  assign new_n14901 = ~new_n14900 & new_n8515;
  assign new_n14902 = n2040 & new_n4138;
  assign new_n14903 = ~new_n14902 & new_n14845;
  assign new_n14904 = ~new_n4643 & ~new_n9302;
  assign new_n14905 = ~new_n9092 & new_n4150;
  assign new_n14906 = ~new_n14904 & ~new_n14905;
  assign new_n14907 = new_n14903 & new_n14906;
  assign new_n14908 = ~new_n14907 & new_n8515;
  assign new_n14909 = n2039 & new_n4138;
  assign new_n14910 = ~new_n14909 & new_n14845;
  assign new_n14911 = ~new_n4667 & ~new_n9302;
  assign new_n14912 = ~new_n9882 & new_n4150;
  assign new_n14913 = ~new_n14911 & ~new_n14912;
  assign new_n14914 = new_n14910 & new_n14913;
  assign new_n14915 = ~new_n14914 & new_n8515;
  assign new_n14916 = n2038 & new_n4138;
  assign new_n14917 = ~new_n14916 & new_n14845;
  assign new_n14918 = ~new_n4595 & ~new_n9302;
  assign new_n14919 = ~new_n10663 & new_n4150;
  assign new_n14920 = ~new_n14918 & ~new_n14919;
  assign new_n14921 = new_n14917 & new_n14920;
  assign new_n14922 = ~new_n14921 & new_n8515;
  assign new_n14923 = n2037 & new_n4138;
  assign new_n14924 = ~new_n14923 & new_n14845;
  assign new_n14925 = ~new_n4620 & ~new_n9302;
  assign new_n14926 = ~new_n11442 & new_n4150;
  assign new_n14927 = ~new_n14925 & ~new_n14926;
  assign new_n14928 = new_n14924 & new_n14927;
  assign new_n14929 = ~new_n14928 & new_n8515;
  assign new_n14930 = n2036 & new_n4138;
  assign new_n14931 = ~new_n14930 & new_n14845;
  assign new_n14932 = ~new_n4527 & ~new_n9302;
  assign new_n14933 = ~new_n12220 & new_n4150;
  assign new_n14934 = ~new_n14932 & ~new_n14933;
  assign new_n14935 = new_n14931 & new_n14934;
  assign new_n14936 = ~new_n14935 & new_n8515;
  assign new_n14937 = n2035 & new_n4138;
  assign new_n14938 = ~new_n14937 & new_n14845;
  assign new_n14939 = ~new_n4565 & ~new_n9302;
  assign new_n14940 = ~new_n12998 & new_n4150;
  assign new_n14941 = ~new_n14939 & ~new_n14940;
  assign new_n14942 = new_n14938 & new_n14941;
  assign new_n14943 = ~new_n14942 & new_n8515;
  assign new_n14944 = n2034 & new_n4138;
  assign new_n14945 = ~new_n14944 & new_n14845;
  assign new_n14946 = ~new_n4401 & ~new_n9302;
  assign new_n14947 = ~new_n13776 & new_n4150;
  assign new_n14948 = ~new_n14946 & ~new_n14947;
  assign new_n14949 = new_n14945 & new_n14948;
  assign new_n14950 = ~new_n14949 & new_n8515;
  assign new_n14951 = n2033 & new_n4138;
  assign new_n14952 = ~new_n14951 & new_n14845;
  assign new_n14953 = ~new_n4479 & ~new_n9302;
  assign new_n14954 = ~new_n14554 & new_n4150;
  assign new_n14955 = ~new_n14953 & ~new_n14954;
  assign new_n14956 = new_n14952 & new_n14955;
  assign new_n14957 = ~new_n14956 & new_n8515;
  assign new_n14958 = ~new_n8512 & new_n8490;
  assign new_n14959 = new_n14958 ^ new_n8490;
  assign new_n14960 = ~new_n8449 & new_n14959;
  assign new_n14961 = ~new_n9310 & new_n14960;
  assign new_n14962 = ~new_n10088 & new_n14960;
  assign new_n14963 = ~new_n10870 & new_n14960;
  assign new_n14964 = ~new_n11648 & new_n14960;
  assign new_n14965 = ~new_n12426 & new_n14960;
  assign new_n14966 = ~new_n13204 & new_n14960;
  assign new_n14967 = ~new_n13982 & new_n14960;
  assign new_n14968 = ~new_n14760 & new_n14960;
  assign new_n14969 = ~new_n14771 & new_n14960;
  assign new_n14970 = ~new_n14781 & new_n14960;
  assign new_n14971 = ~new_n14791 & new_n14960;
  assign new_n14972 = ~new_n14801 & new_n14960;
  assign new_n14973 = ~new_n14811 & new_n14960;
  assign new_n14974 = ~new_n14821 & new_n14960;
  assign new_n14975 = ~new_n14831 & new_n14960;
  assign new_n14976 = ~new_n14841 & new_n14960;
  assign new_n14977 = ~new_n14851 & new_n14960;
  assign new_n14978 = ~new_n14858 & new_n14960;
  assign new_n14979 = ~new_n14865 & new_n14960;
  assign new_n14980 = ~new_n14872 & new_n14960;
  assign new_n14981 = ~new_n14879 & new_n14960;
  assign new_n14982 = ~new_n14886 & new_n14960;
  assign new_n14983 = ~new_n14893 & new_n14960;
  assign new_n14984 = ~new_n14900 & new_n14960;
  assign new_n14985 = ~new_n14907 & new_n14960;
  assign new_n14986 = ~new_n14914 & new_n14960;
  assign new_n14987 = ~new_n14921 & new_n14960;
  assign new_n14988 = ~new_n14928 & new_n14960;
  assign new_n14989 = ~new_n14935 & new_n14960;
  assign new_n14990 = ~new_n14942 & new_n14960;
  assign new_n14991 = ~new_n14949 & new_n14960;
  assign new_n14992 = ~new_n14956 & new_n14960;
  assign new_n14993 = ~new_n8491 & ~new_n8512;
  assign new_n14994 = new_n14993 ^ new_n8491;
  assign new_n14995 = ~new_n8449 & ~new_n14994;
  assign new_n14996 = ~new_n9310 & new_n14995;
  assign new_n14997 = ~new_n10088 & new_n14995;
  assign new_n14998 = ~new_n10870 & new_n14995;
  assign new_n14999 = ~new_n11648 & new_n14995;
  assign new_n15000 = ~new_n12426 & new_n14995;
  assign new_n15001 = ~new_n13204 & new_n14995;
  assign new_n15002 = ~new_n13982 & new_n14995;
  assign new_n15003 = ~new_n14760 & new_n14995;
  assign new_n15004 = ~new_n14771 & new_n14995;
  assign new_n15005 = ~new_n14781 & new_n14995;
  assign new_n15006 = ~new_n14791 & new_n14995;
  assign new_n15007 = ~new_n14801 & new_n14995;
  assign new_n15008 = ~new_n14811 & new_n14995;
  assign new_n15009 = ~new_n14821 & new_n14995;
  assign new_n15010 = ~new_n14831 & new_n14995;
  assign new_n15011 = ~new_n14841 & new_n14995;
  assign new_n15012 = ~new_n14851 & new_n14995;
  assign new_n15013 = ~new_n14858 & new_n14995;
  assign new_n15014 = ~new_n14865 & new_n14995;
  assign new_n15015 = ~new_n14872 & new_n14995;
  assign new_n15016 = ~new_n14879 & new_n14995;
  assign new_n15017 = ~new_n14886 & new_n14995;
  assign new_n15018 = ~new_n14893 & new_n14995;
  assign new_n15019 = ~new_n14900 & new_n14995;
  assign new_n15020 = ~new_n14907 & new_n14995;
  assign new_n15021 = ~new_n14914 & new_n14995;
  assign new_n15022 = ~new_n14921 & new_n14995;
  assign new_n15023 = ~new_n14928 & new_n14995;
  assign new_n15024 = ~new_n14935 & new_n14995;
  assign new_n15025 = ~new_n14942 & new_n14995;
  assign new_n15026 = ~new_n14949 & new_n14995;
  assign new_n15027 = ~new_n14956 & new_n14995;
  assign new_n15028 = new_n8489 & new_n8512;
  assign new_n15029 = new_n15028 ^ new_n8489;
  assign new_n15030 = ~new_n8449 & new_n15029;
  assign new_n15031 = ~new_n9310 & new_n15030;
  assign new_n15032 = ~new_n10088 & new_n15030;
  assign new_n15033 = ~new_n10870 & new_n15030;
  assign new_n15034 = ~new_n11648 & new_n15030;
  assign new_n15035 = ~new_n12426 & new_n15030;
  assign new_n15036 = ~new_n13204 & new_n15030;
  assign new_n15037 = ~new_n13982 & new_n15030;
  assign new_n15038 = ~new_n14760 & new_n15030;
  assign new_n15039 = ~new_n14771 & new_n15030;
  assign new_n15040 = ~new_n14781 & new_n15030;
  assign new_n15041 = ~new_n14791 & new_n15030;
  assign new_n15042 = ~new_n14801 & new_n15030;
  assign new_n15043 = ~new_n14811 & new_n15030;
  assign new_n15044 = ~new_n14821 & new_n15030;
  assign new_n15045 = ~new_n14831 & new_n15030;
  assign new_n15046 = ~new_n14841 & new_n15030;
  assign new_n15047 = ~new_n14851 & new_n15030;
  assign new_n15048 = ~new_n14858 & new_n15030;
  assign new_n15049 = ~new_n14865 & new_n15030;
  assign new_n15050 = ~new_n14872 & new_n15030;
  assign new_n15051 = ~new_n14879 & new_n15030;
  assign new_n15052 = ~new_n14886 & new_n15030;
  assign new_n15053 = ~new_n14893 & new_n15030;
  assign new_n15054 = ~new_n14900 & new_n15030;
  assign new_n15055 = ~new_n14907 & new_n15030;
  assign new_n15056 = ~new_n14914 & new_n15030;
  assign new_n15057 = ~new_n14921 & new_n15030;
  assign new_n15058 = ~new_n14928 & new_n15030;
  assign new_n15059 = ~new_n14935 & new_n15030;
  assign new_n15060 = ~new_n14942 & new_n15030;
  assign new_n15061 = ~new_n14949 & new_n15030;
  assign new_n15062 = ~new_n14956 & new_n15030;
  assign new_n15063 = ~new_n8449 & new_n8513;
  assign new_n15064 = ~new_n9310 & new_n15063;
  assign new_n15065 = ~new_n10088 & new_n15063;
  assign new_n15066 = ~new_n10870 & new_n15063;
  assign new_n15067 = ~new_n11648 & new_n15063;
  assign new_n15068 = ~new_n12426 & new_n15063;
  assign new_n15069 = ~new_n13204 & new_n15063;
  assign new_n15070 = ~new_n13982 & new_n15063;
  assign new_n15071 = ~new_n14760 & new_n15063;
  assign new_n15072 = ~new_n14771 & new_n15063;
  assign new_n15073 = ~new_n14781 & new_n15063;
  assign new_n15074 = ~new_n14791 & new_n15063;
  assign new_n15075 = ~new_n14801 & new_n15063;
  assign new_n15076 = ~new_n14811 & new_n15063;
  assign new_n15077 = ~new_n14821 & new_n15063;
  assign new_n15078 = ~new_n14831 & new_n15063;
  assign new_n15079 = ~new_n14841 & new_n15063;
  assign new_n15080 = ~new_n14851 & new_n15063;
  assign new_n15081 = ~new_n14858 & new_n15063;
  assign new_n15082 = ~new_n14865 & new_n15063;
  assign new_n15083 = ~new_n14872 & new_n15063;
  assign new_n15084 = ~new_n14879 & new_n15063;
  assign new_n15085 = ~new_n14886 & new_n15063;
  assign new_n15086 = ~new_n14893 & new_n15063;
  assign new_n15087 = ~new_n14900 & new_n15063;
  assign new_n15088 = ~new_n14907 & new_n15063;
  assign new_n15089 = ~new_n14914 & new_n15063;
  assign new_n15090 = ~new_n14921 & new_n15063;
  assign new_n15091 = ~new_n14928 & new_n15063;
  assign new_n15092 = ~new_n14935 & new_n15063;
  assign new_n15093 = ~new_n14942 & new_n15063;
  assign new_n15094 = ~new_n14949 & new_n15063;
  assign new_n15095 = ~new_n14956 & new_n15063;
  assign new_n15096 = ~new_n8449 & new_n14958;
  assign new_n15097 = ~new_n9310 & new_n15096;
  assign new_n15098 = ~new_n10088 & new_n15096;
  assign new_n15099 = ~new_n10870 & new_n15096;
  assign new_n15100 = ~new_n11648 & new_n15096;
  assign new_n15101 = ~new_n12426 & new_n15096;
  assign new_n15102 = ~new_n13204 & new_n15096;
  assign new_n15103 = ~new_n13982 & new_n15096;
  assign new_n15104 = ~new_n14760 & new_n15096;
  assign new_n15105 = ~new_n14771 & new_n15096;
  assign new_n15106 = ~new_n14781 & new_n15096;
  assign new_n15107 = ~new_n14791 & new_n15096;
  assign new_n15108 = ~new_n14801 & new_n15096;
  assign new_n15109 = ~new_n14811 & new_n15096;
  assign new_n15110 = ~new_n14821 & new_n15096;
  assign new_n15111 = ~new_n14831 & new_n15096;
  assign new_n15112 = ~new_n14841 & new_n15096;
  assign new_n15113 = ~new_n14851 & new_n15096;
  assign new_n15114 = ~new_n14858 & new_n15096;
  assign new_n15115 = ~new_n14865 & new_n15096;
  assign new_n15116 = ~new_n14872 & new_n15096;
  assign new_n15117 = ~new_n14879 & new_n15096;
  assign new_n15118 = ~new_n14886 & new_n15096;
  assign new_n15119 = ~new_n14893 & new_n15096;
  assign new_n15120 = ~new_n14900 & new_n15096;
  assign new_n15121 = ~new_n14907 & new_n15096;
  assign new_n15122 = ~new_n14914 & new_n15096;
  assign new_n15123 = ~new_n14921 & new_n15096;
  assign new_n15124 = ~new_n14928 & new_n15096;
  assign new_n15125 = ~new_n14935 & new_n15096;
  assign new_n15126 = ~new_n14942 & new_n15096;
  assign new_n15127 = ~new_n14949 & new_n15096;
  assign new_n15128 = ~new_n14956 & new_n15096;
  assign new_n15129 = ~new_n8449 & new_n14993;
  assign new_n15130 = ~new_n9310 & new_n15129;
  assign new_n15131 = ~new_n10088 & new_n15129;
  assign new_n15132 = ~new_n10870 & new_n15129;
  assign new_n15133 = ~new_n11648 & new_n15129;
  assign new_n15134 = ~new_n12426 & new_n15129;
  assign new_n15135 = ~new_n13204 & new_n15129;
  assign new_n15136 = ~new_n13982 & new_n15129;
  assign new_n15137 = ~new_n14760 & new_n15129;
  assign new_n15138 = ~new_n14771 & new_n15129;
  assign new_n15139 = ~new_n14781 & new_n15129;
  assign new_n15140 = ~new_n14791 & new_n15129;
  assign new_n15141 = ~new_n14801 & new_n15129;
  assign new_n15142 = ~new_n14811 & new_n15129;
  assign new_n15143 = ~new_n14821 & new_n15129;
  assign new_n15144 = ~new_n14831 & new_n15129;
  assign new_n15145 = ~new_n14841 & new_n15129;
  assign new_n15146 = ~new_n14851 & new_n15129;
  assign new_n15147 = ~new_n14858 & new_n15129;
  assign new_n15148 = ~new_n14865 & new_n15129;
  assign new_n15149 = ~new_n14872 & new_n15129;
  assign new_n15150 = ~new_n14879 & new_n15129;
  assign new_n15151 = ~new_n14886 & new_n15129;
  assign new_n15152 = ~new_n14893 & new_n15129;
  assign new_n15153 = ~new_n14900 & new_n15129;
  assign new_n15154 = ~new_n14907 & new_n15129;
  assign new_n15155 = ~new_n14914 & new_n15129;
  assign new_n15156 = ~new_n14921 & new_n15129;
  assign new_n15157 = ~new_n14928 & new_n15129;
  assign new_n15158 = ~new_n14935 & new_n15129;
  assign new_n15159 = ~new_n14942 & new_n15129;
  assign new_n15160 = ~new_n14949 & new_n15129;
  assign new_n15161 = ~new_n14956 & new_n15129;
  assign new_n15162 = new_n8447 ^ new_n8427;
  assign new_n15163 = ~new_n15162 & new_n15028;
  assign new_n15164 = ~new_n9310 & new_n15163;
  assign new_n15165 = ~new_n10088 & new_n15163;
  assign new_n15166 = ~new_n10870 & new_n15163;
  assign new_n15167 = ~new_n11648 & new_n15163;
  assign new_n15168 = ~new_n12426 & new_n15163;
  assign new_n15169 = ~new_n13204 & new_n15163;
  assign new_n15170 = ~new_n13982 & new_n15163;
  assign new_n15171 = ~new_n14760 & new_n15163;
  assign new_n15172 = ~new_n14771 & new_n15163;
  assign new_n15173 = ~new_n14781 & new_n15163;
  assign new_n15174 = ~new_n14791 & new_n15163;
  assign new_n15175 = ~new_n14801 & new_n15163;
  assign new_n15176 = ~new_n14811 & new_n15163;
  assign new_n15177 = ~new_n14821 & new_n15163;
  assign new_n15178 = ~new_n14831 & new_n15163;
  assign new_n15179 = ~new_n14841 & new_n15163;
  assign new_n15180 = ~new_n14851 & new_n15163;
  assign new_n15181 = ~new_n14858 & new_n15163;
  assign new_n15182 = ~new_n14865 & new_n15163;
  assign new_n15183 = ~new_n14872 & new_n15163;
  assign new_n15184 = ~new_n14879 & new_n15163;
  assign new_n15185 = ~new_n14886 & new_n15163;
  assign new_n15186 = ~new_n14893 & new_n15163;
  assign new_n15187 = ~new_n14900 & new_n15163;
  assign new_n15188 = ~new_n14907 & new_n15163;
  assign new_n15189 = ~new_n14914 & new_n15163;
  assign new_n15190 = ~new_n14921 & new_n15163;
  assign new_n15191 = ~new_n14928 & new_n15163;
  assign new_n15192 = ~new_n14935 & new_n15163;
  assign new_n15193 = ~new_n14942 & new_n15163;
  assign new_n15194 = ~new_n14949 & new_n15163;
  assign new_n15195 = ~new_n14956 & new_n15163;
  assign new_n15196 = ~new_n15162 & new_n8514;
  assign new_n15197 = ~new_n9310 & new_n15196;
  assign new_n15198 = ~new_n10088 & new_n15196;
  assign new_n15199 = ~new_n10870 & new_n15196;
  assign new_n15200 = ~new_n11648 & new_n15196;
  assign new_n15201 = ~new_n12426 & new_n15196;
  assign new_n15202 = ~new_n13204 & new_n15196;
  assign new_n15203 = ~new_n13982 & new_n15196;
  assign new_n15204 = ~new_n14760 & new_n15196;
  assign new_n15205 = ~new_n14771 & new_n15196;
  assign new_n15206 = ~new_n14781 & new_n15196;
  assign new_n15207 = ~new_n14791 & new_n15196;
  assign new_n15208 = ~new_n14801 & new_n15196;
  assign new_n15209 = ~new_n14811 & new_n15196;
  assign new_n15210 = ~new_n14821 & new_n15196;
  assign new_n15211 = ~new_n14831 & new_n15196;
  assign new_n15212 = ~new_n14841 & new_n15196;
  assign new_n15213 = ~new_n14851 & new_n15196;
  assign new_n15214 = ~new_n14858 & new_n15196;
  assign new_n15215 = ~new_n14865 & new_n15196;
  assign new_n15216 = ~new_n14872 & new_n15196;
  assign new_n15217 = ~new_n14879 & new_n15196;
  assign new_n15218 = ~new_n14886 & new_n15196;
  assign new_n15219 = ~new_n14893 & new_n15196;
  assign new_n15220 = ~new_n14900 & new_n15196;
  assign new_n15221 = ~new_n14907 & new_n15196;
  assign new_n15222 = ~new_n14914 & new_n15196;
  assign new_n15223 = ~new_n14921 & new_n15196;
  assign new_n15224 = ~new_n14928 & new_n15196;
  assign new_n15225 = ~new_n14935 & new_n15196;
  assign new_n15226 = ~new_n14942 & new_n15196;
  assign new_n15227 = ~new_n14949 & new_n15196;
  assign new_n15228 = ~new_n14956 & new_n15196;
  assign new_n15229 = ~new_n15162 & new_n14959;
  assign new_n15230 = ~new_n9310 & new_n15229;
  assign new_n15231 = ~new_n10088 & new_n15229;
  assign new_n15232 = ~new_n10870 & new_n15229;
  assign new_n15233 = ~new_n11648 & new_n15229;
  assign new_n15234 = ~new_n12426 & new_n15229;
  assign new_n15235 = ~new_n13204 & new_n15229;
  assign new_n15236 = ~new_n13982 & new_n15229;
  assign new_n15237 = ~new_n14760 & new_n15229;
  assign new_n15238 = ~new_n14771 & new_n15229;
  assign new_n15239 = ~new_n14781 & new_n15229;
  assign new_n15240 = ~new_n14791 & new_n15229;
  assign new_n15241 = ~new_n14801 & new_n15229;
  assign new_n15242 = ~new_n14811 & new_n15229;
  assign new_n15243 = ~new_n14821 & new_n15229;
  assign new_n15244 = ~new_n14831 & new_n15229;
  assign new_n15245 = ~new_n14841 & new_n15229;
  assign new_n15246 = ~new_n14851 & new_n15229;
  assign new_n15247 = ~new_n14858 & new_n15229;
  assign new_n15248 = ~new_n14865 & new_n15229;
  assign new_n15249 = ~new_n14872 & new_n15229;
  assign new_n15250 = ~new_n14879 & new_n15229;
  assign new_n15251 = ~new_n14886 & new_n15229;
  assign new_n15252 = ~new_n14893 & new_n15229;
  assign new_n15253 = ~new_n14900 & new_n15229;
  assign new_n15254 = ~new_n14907 & new_n15229;
  assign new_n15255 = ~new_n14914 & new_n15229;
  assign new_n15256 = ~new_n14921 & new_n15229;
  assign new_n15257 = ~new_n14928 & new_n15229;
  assign new_n15258 = ~new_n14935 & new_n15229;
  assign new_n15259 = ~new_n14942 & new_n15229;
  assign new_n15260 = ~new_n14949 & new_n15229;
  assign new_n15261 = ~new_n14956 & new_n15229;
  assign new_n15262 = ~new_n14994 & ~new_n15162;
  assign new_n15263 = ~new_n9310 & new_n15262;
  assign new_n15264 = ~new_n10088 & new_n15262;
  assign new_n15265 = ~new_n10870 & new_n15262;
  assign new_n15266 = ~new_n11648 & new_n15262;
  assign new_n15267 = ~new_n12426 & new_n15262;
  assign new_n15268 = ~new_n13204 & new_n15262;
  assign new_n15269 = ~new_n13982 & new_n15262;
  assign new_n15270 = ~new_n14760 & new_n15262;
  assign new_n15271 = ~new_n14771 & new_n15262;
  assign new_n15272 = ~new_n14781 & new_n15262;
  assign new_n15273 = ~new_n14791 & new_n15262;
  assign new_n15274 = ~new_n14801 & new_n15262;
  assign new_n15275 = ~new_n14811 & new_n15262;
  assign new_n15276 = ~new_n14821 & new_n15262;
  assign new_n15277 = ~new_n14831 & new_n15262;
  assign new_n15278 = ~new_n14841 & new_n15262;
  assign new_n15279 = ~new_n14851 & new_n15262;
  assign new_n15280 = ~new_n14858 & new_n15262;
  assign new_n15281 = ~new_n14865 & new_n15262;
  assign new_n15282 = ~new_n14872 & new_n15262;
  assign new_n15283 = ~new_n14879 & new_n15262;
  assign new_n15284 = ~new_n14886 & new_n15262;
  assign new_n15285 = ~new_n14893 & new_n15262;
  assign new_n15286 = ~new_n14900 & new_n15262;
  assign new_n15287 = ~new_n14907 & new_n15262;
  assign new_n15288 = ~new_n14914 & new_n15262;
  assign new_n15289 = ~new_n14921 & new_n15262;
  assign new_n15290 = ~new_n14928 & new_n15262;
  assign new_n15291 = ~new_n14935 & new_n15262;
  assign new_n15292 = ~new_n14942 & new_n15262;
  assign new_n15293 = ~new_n14949 & new_n15262;
  assign new_n15294 = ~new_n14956 & new_n15262;
  assign new_n15295 = ~new_n15162 & new_n15029;
  assign new_n15296 = ~new_n9310 & new_n15295;
  assign new_n15297 = ~new_n10088 & new_n15295;
  assign new_n15298 = ~new_n10870 & new_n15295;
  assign new_n15299 = ~new_n11648 & new_n15295;
  assign new_n15300 = ~new_n12426 & new_n15295;
  assign new_n15301 = ~new_n13204 & new_n15295;
  assign new_n15302 = ~new_n13982 & new_n15295;
  assign new_n15303 = ~new_n14760 & new_n15295;
  assign new_n15304 = ~new_n14771 & new_n15295;
  assign new_n15305 = ~new_n14781 & new_n15295;
  assign new_n15306 = ~new_n14791 & new_n15295;
  assign new_n15307 = ~new_n14801 & new_n15295;
  assign new_n15308 = ~new_n14811 & new_n15295;
  assign new_n15309 = ~new_n14821 & new_n15295;
  assign new_n15310 = ~new_n14831 & new_n15295;
  assign new_n15311 = ~new_n14841 & new_n15295;
  assign new_n15312 = ~new_n14851 & new_n15295;
  assign new_n15313 = ~new_n14858 & new_n15295;
  assign new_n15314 = ~new_n14865 & new_n15295;
  assign new_n15315 = ~new_n14872 & new_n15295;
  assign new_n15316 = ~new_n14879 & new_n15295;
  assign new_n15317 = ~new_n14886 & new_n15295;
  assign new_n15318 = ~new_n14893 & new_n15295;
  assign new_n15319 = ~new_n14900 & new_n15295;
  assign new_n15320 = ~new_n14907 & new_n15295;
  assign new_n15321 = ~new_n14914 & new_n15295;
  assign new_n15322 = ~new_n14921 & new_n15295;
  assign new_n15323 = ~new_n14928 & new_n15295;
  assign new_n15324 = ~new_n14935 & new_n15295;
  assign new_n15325 = ~new_n14942 & new_n15295;
  assign new_n15326 = ~new_n14949 & new_n15295;
  assign new_n15327 = ~new_n14956 & new_n15295;
  assign new_n15328 = ~new_n15162 & new_n8513;
  assign new_n15329 = ~new_n9310 & new_n15328;
  assign new_n15330 = ~new_n10088 & new_n15328;
  assign new_n15331 = ~new_n10870 & new_n15328;
  assign new_n15332 = ~new_n11648 & new_n15328;
  assign new_n15333 = ~new_n12426 & new_n15328;
  assign new_n15334 = ~new_n13204 & new_n15328;
  assign new_n15335 = ~new_n13982 & new_n15328;
  assign new_n15336 = ~new_n14760 & new_n15328;
  assign new_n15337 = ~new_n14771 & new_n15328;
  assign new_n15338 = ~new_n14781 & new_n15328;
  assign new_n15339 = ~new_n14791 & new_n15328;
  assign new_n15340 = ~new_n14801 & new_n15328;
  assign new_n15341 = ~new_n14811 & new_n15328;
  assign new_n15342 = ~new_n14821 & new_n15328;
  assign new_n15343 = ~new_n14831 & new_n15328;
  assign new_n15344 = ~new_n14841 & new_n15328;
  assign new_n15345 = ~new_n14851 & new_n15328;
  assign new_n15346 = ~new_n14858 & new_n15328;
  assign new_n15347 = ~new_n14865 & new_n15328;
  assign new_n15348 = ~new_n14872 & new_n15328;
  assign new_n15349 = ~new_n14879 & new_n15328;
  assign new_n15350 = ~new_n14886 & new_n15328;
  assign new_n15351 = ~new_n14893 & new_n15328;
  assign new_n15352 = ~new_n14900 & new_n15328;
  assign new_n15353 = ~new_n14907 & new_n15328;
  assign new_n15354 = ~new_n14914 & new_n15328;
  assign new_n15355 = ~new_n14921 & new_n15328;
  assign new_n15356 = ~new_n14928 & new_n15328;
  assign new_n15357 = ~new_n14935 & new_n15328;
  assign new_n15358 = ~new_n14942 & new_n15328;
  assign new_n15359 = ~new_n14949 & new_n15328;
  assign new_n15360 = ~new_n14956 & new_n15328;
  assign new_n15361 = ~new_n15162 & new_n14958;
  assign new_n15362 = ~new_n9310 & new_n15361;
  assign new_n15363 = ~new_n10088 & new_n15361;
  assign new_n15364 = ~new_n10870 & new_n15361;
  assign new_n15365 = ~new_n11648 & new_n15361;
  assign new_n15366 = ~new_n12426 & new_n15361;
  assign new_n15367 = ~new_n13204 & new_n15361;
  assign new_n15368 = ~new_n13982 & new_n15361;
  assign new_n15369 = ~new_n14760 & new_n15361;
  assign new_n15370 = ~new_n14771 & new_n15361;
  assign new_n15371 = ~new_n14781 & new_n15361;
  assign new_n15372 = ~new_n14791 & new_n15361;
  assign new_n15373 = ~new_n14801 & new_n15361;
  assign new_n15374 = ~new_n14811 & new_n15361;
  assign new_n15375 = ~new_n14821 & new_n15361;
  assign new_n15376 = ~new_n14831 & new_n15361;
  assign new_n15377 = ~new_n14841 & new_n15361;
  assign new_n15378 = ~new_n14851 & new_n15361;
  assign new_n15379 = ~new_n14858 & new_n15361;
  assign new_n15380 = ~new_n14865 & new_n15361;
  assign new_n15381 = ~new_n14872 & new_n15361;
  assign new_n15382 = ~new_n14879 & new_n15361;
  assign new_n15383 = ~new_n14886 & new_n15361;
  assign new_n15384 = ~new_n14893 & new_n15361;
  assign new_n15385 = ~new_n14900 & new_n15361;
  assign new_n15386 = ~new_n14907 & new_n15361;
  assign new_n15387 = ~new_n14914 & new_n15361;
  assign new_n15388 = ~new_n14921 & new_n15361;
  assign new_n15389 = ~new_n14928 & new_n15361;
  assign new_n15390 = ~new_n14935 & new_n15361;
  assign new_n15391 = ~new_n14942 & new_n15361;
  assign new_n15392 = ~new_n14949 & new_n15361;
  assign new_n15393 = ~new_n14956 & new_n15361;
  assign new_n15394 = ~new_n15162 & new_n14993;
  assign new_n15395 = ~new_n9310 & new_n15394;
  assign new_n15396 = ~new_n10088 & new_n15394;
  assign new_n15397 = ~new_n10870 & new_n15394;
  assign new_n15398 = ~new_n11648 & new_n15394;
  assign new_n15399 = ~new_n12426 & new_n15394;
  assign new_n15400 = ~new_n13204 & new_n15394;
  assign new_n15401 = ~new_n13982 & new_n15394;
  assign new_n15402 = ~new_n14760 & new_n15394;
  assign new_n15403 = ~new_n14771 & new_n15394;
  assign new_n15404 = ~new_n14781 & new_n15394;
  assign new_n15405 = ~new_n14791 & new_n15394;
  assign new_n15406 = ~new_n14801 & new_n15394;
  assign new_n15407 = ~new_n14811 & new_n15394;
  assign new_n15408 = ~new_n14821 & new_n15394;
  assign new_n15409 = ~new_n14831 & new_n15394;
  assign new_n15410 = ~new_n14841 & new_n15394;
  assign new_n15411 = ~new_n14851 & new_n15394;
  assign new_n15412 = ~new_n14858 & new_n15394;
  assign new_n15413 = ~new_n14865 & new_n15394;
  assign new_n15414 = ~new_n14872 & new_n15394;
  assign new_n15415 = ~new_n14879 & new_n15394;
  assign new_n15416 = ~new_n14886 & new_n15394;
  assign new_n15417 = ~new_n14893 & new_n15394;
  assign new_n15418 = ~new_n14900 & new_n15394;
  assign new_n15419 = ~new_n14907 & new_n15394;
  assign new_n15420 = ~new_n14914 & new_n15394;
  assign new_n15421 = ~new_n14921 & new_n15394;
  assign new_n15422 = ~new_n14928 & new_n15394;
  assign new_n15423 = ~new_n14935 & new_n15394;
  assign new_n15424 = ~new_n14942 & new_n15394;
  assign new_n15425 = ~new_n14949 & new_n15394;
  assign new_n15426 = ~new_n14956 & new_n15394;
  assign new_n15427 = ~new_n8448 & new_n15028;
  assign new_n15428 = ~new_n9310 & new_n15427;
  assign new_n15429 = ~new_n10088 & new_n15427;
  assign new_n15430 = ~new_n10870 & new_n15427;
  assign new_n15431 = ~new_n11648 & new_n15427;
  assign new_n15432 = ~new_n12426 & new_n15427;
  assign new_n15433 = ~new_n13204 & new_n15427;
  assign new_n15434 = ~new_n13982 & new_n15427;
  assign new_n15435 = ~new_n14760 & new_n15427;
  assign new_n15436 = ~new_n14771 & new_n15427;
  assign new_n15437 = ~new_n14781 & new_n15427;
  assign new_n15438 = ~new_n14791 & new_n15427;
  assign new_n15439 = ~new_n14801 & new_n15427;
  assign new_n15440 = ~new_n14811 & new_n15427;
  assign new_n15441 = ~new_n14821 & new_n15427;
  assign new_n15442 = ~new_n14831 & new_n15427;
  assign new_n15443 = ~new_n14841 & new_n15427;
  assign new_n15444 = ~new_n14851 & new_n15427;
  assign new_n15445 = ~new_n14858 & new_n15427;
  assign new_n15446 = ~new_n14865 & new_n15427;
  assign new_n15447 = ~new_n14872 & new_n15427;
  assign new_n15448 = ~new_n14879 & new_n15427;
  assign new_n15449 = ~new_n14886 & new_n15427;
  assign new_n15450 = ~new_n14893 & new_n15427;
  assign new_n15451 = ~new_n14900 & new_n15427;
  assign new_n15452 = ~new_n14907 & new_n15427;
  assign new_n15453 = ~new_n14914 & new_n15427;
  assign new_n15454 = ~new_n14921 & new_n15427;
  assign new_n15455 = ~new_n14928 & new_n15427;
  assign new_n15456 = ~new_n14935 & new_n15427;
  assign new_n15457 = ~new_n14942 & new_n15427;
  assign new_n15458 = ~new_n14949 & new_n15427;
  assign new_n15459 = ~new_n14956 & new_n15427;
  assign new_n15460 = ~new_n8448 & new_n8514;
  assign new_n15461 = ~new_n9310 & new_n15460;
  assign new_n15462 = ~new_n10088 & new_n15460;
  assign new_n15463 = ~new_n10870 & new_n15460;
  assign new_n15464 = ~new_n11648 & new_n15460;
  assign new_n15465 = ~new_n12426 & new_n15460;
  assign new_n15466 = ~new_n13204 & new_n15460;
  assign new_n15467 = ~new_n13982 & new_n15460;
  assign new_n15468 = ~new_n14760 & new_n15460;
  assign new_n15469 = ~new_n14771 & new_n15460;
  assign new_n15470 = ~new_n14781 & new_n15460;
  assign new_n15471 = ~new_n14791 & new_n15460;
  assign new_n15472 = ~new_n14801 & new_n15460;
  assign new_n15473 = ~new_n14811 & new_n15460;
  assign new_n15474 = ~new_n14821 & new_n15460;
  assign new_n15475 = ~new_n14831 & new_n15460;
  assign new_n15476 = ~new_n14841 & new_n15460;
  assign new_n15477 = ~new_n14851 & new_n15460;
  assign new_n15478 = ~new_n14858 & new_n15460;
  assign new_n15479 = ~new_n14865 & new_n15460;
  assign new_n15480 = ~new_n14872 & new_n15460;
  assign new_n15481 = ~new_n14879 & new_n15460;
  assign new_n15482 = ~new_n14886 & new_n15460;
  assign new_n15483 = ~new_n14893 & new_n15460;
  assign new_n15484 = ~new_n14900 & new_n15460;
  assign new_n15485 = ~new_n14907 & new_n15460;
  assign new_n15486 = ~new_n14914 & new_n15460;
  assign new_n15487 = ~new_n14921 & new_n15460;
  assign new_n15488 = ~new_n14928 & new_n15460;
  assign new_n15489 = ~new_n14935 & new_n15460;
  assign new_n15490 = ~new_n14942 & new_n15460;
  assign new_n15491 = ~new_n14949 & new_n15460;
  assign new_n15492 = ~new_n14956 & new_n15460;
  assign new_n15493 = ~new_n8448 & new_n14959;
  assign new_n15494 = ~new_n9310 & new_n15493;
  assign new_n15495 = ~new_n10088 & new_n15493;
  assign new_n15496 = ~new_n10870 & new_n15493;
  assign new_n15497 = ~new_n11648 & new_n15493;
  assign new_n15498 = ~new_n12426 & new_n15493;
  assign new_n15499 = ~new_n13204 & new_n15493;
  assign new_n15500 = ~new_n13982 & new_n15493;
  assign new_n15501 = ~new_n14760 & new_n15493;
  assign new_n15502 = ~new_n14771 & new_n15493;
  assign new_n15503 = ~new_n14781 & new_n15493;
  assign new_n15504 = ~new_n14791 & new_n15493;
  assign new_n15505 = ~new_n14801 & new_n15493;
  assign new_n15506 = ~new_n14811 & new_n15493;
  assign new_n15507 = ~new_n14821 & new_n15493;
  assign new_n15508 = ~new_n14831 & new_n15493;
  assign new_n15509 = ~new_n14841 & new_n15493;
  assign new_n15510 = ~new_n14851 & new_n15493;
  assign new_n15511 = ~new_n14858 & new_n15493;
  assign new_n15512 = ~new_n14865 & new_n15493;
  assign new_n15513 = ~new_n14872 & new_n15493;
  assign new_n15514 = ~new_n14879 & new_n15493;
  assign new_n15515 = ~new_n14886 & new_n15493;
  assign new_n15516 = ~new_n14893 & new_n15493;
  assign new_n15517 = ~new_n14900 & new_n15493;
  assign new_n15518 = ~new_n14907 & new_n15493;
  assign new_n15519 = ~new_n14914 & new_n15493;
  assign new_n15520 = ~new_n14921 & new_n15493;
  assign new_n15521 = ~new_n14928 & new_n15493;
  assign new_n15522 = ~new_n14935 & new_n15493;
  assign new_n15523 = ~new_n14942 & new_n15493;
  assign new_n15524 = ~new_n14949 & new_n15493;
  assign new_n15525 = ~new_n14956 & new_n15493;
  assign new_n15526 = ~new_n8448 & ~new_n14994;
  assign new_n15527 = ~new_n9310 & new_n15526;
  assign new_n15528 = ~new_n10088 & new_n15526;
  assign new_n15529 = ~new_n10870 & new_n15526;
  assign new_n15530 = ~new_n11648 & new_n15526;
  assign new_n15531 = ~new_n12426 & new_n15526;
  assign new_n15532 = ~new_n13204 & new_n15526;
  assign new_n15533 = ~new_n13982 & new_n15526;
  assign new_n15534 = ~new_n14760 & new_n15526;
  assign new_n15535 = ~new_n14771 & new_n15526;
  assign new_n15536 = ~new_n14781 & new_n15526;
  assign new_n15537 = ~new_n14791 & new_n15526;
  assign new_n15538 = ~new_n14801 & new_n15526;
  assign new_n15539 = ~new_n14811 & new_n15526;
  assign new_n15540 = ~new_n14821 & new_n15526;
  assign new_n15541 = ~new_n14831 & new_n15526;
  assign new_n15542 = ~new_n14841 & new_n15526;
  assign new_n15543 = ~new_n14851 & new_n15526;
  assign new_n15544 = ~new_n14858 & new_n15526;
  assign new_n15545 = ~new_n14865 & new_n15526;
  assign new_n15546 = ~new_n14872 & new_n15526;
  assign new_n15547 = ~new_n14879 & new_n15526;
  assign new_n15548 = ~new_n14886 & new_n15526;
  assign new_n15549 = ~new_n14893 & new_n15526;
  assign new_n15550 = ~new_n14900 & new_n15526;
  assign new_n15551 = ~new_n14907 & new_n15526;
  assign new_n15552 = ~new_n14914 & new_n15526;
  assign new_n15553 = ~new_n14921 & new_n15526;
  assign new_n15554 = ~new_n14928 & new_n15526;
  assign new_n15555 = ~new_n14935 & new_n15526;
  assign new_n15556 = ~new_n14942 & new_n15526;
  assign new_n15557 = ~new_n14949 & new_n15526;
  assign new_n15558 = ~new_n14956 & new_n15526;
  assign new_n15559 = ~new_n8448 & new_n15029;
  assign new_n15560 = ~new_n9310 & new_n15559;
  assign new_n15561 = ~new_n10088 & new_n15559;
  assign new_n15562 = ~new_n10870 & new_n15559;
  assign new_n15563 = ~new_n11648 & new_n15559;
  assign new_n15564 = ~new_n12426 & new_n15559;
  assign new_n15565 = ~new_n13204 & new_n15559;
  assign new_n15566 = ~new_n13982 & new_n15559;
  assign new_n15567 = ~new_n14760 & new_n15559;
  assign new_n15568 = ~new_n14771 & new_n15559;
  assign new_n15569 = ~new_n14781 & new_n15559;
  assign new_n15570 = ~new_n14791 & new_n15559;
  assign new_n15571 = ~new_n14801 & new_n15559;
  assign new_n15572 = ~new_n14811 & new_n15559;
  assign new_n15573 = ~new_n14821 & new_n15559;
  assign new_n15574 = ~new_n14831 & new_n15559;
  assign new_n15575 = ~new_n14841 & new_n15559;
  assign new_n15576 = ~new_n14851 & new_n15559;
  assign new_n15577 = ~new_n14858 & new_n15559;
  assign new_n15578 = ~new_n14865 & new_n15559;
  assign new_n15579 = ~new_n14872 & new_n15559;
  assign new_n15580 = ~new_n14879 & new_n15559;
  assign new_n15581 = ~new_n14886 & new_n15559;
  assign new_n15582 = ~new_n14893 & new_n15559;
  assign new_n15583 = ~new_n14900 & new_n15559;
  assign new_n15584 = ~new_n14907 & new_n15559;
  assign new_n15585 = ~new_n14914 & new_n15559;
  assign new_n15586 = ~new_n14921 & new_n15559;
  assign new_n15587 = ~new_n14928 & new_n15559;
  assign new_n15588 = ~new_n14935 & new_n15559;
  assign new_n15589 = ~new_n14942 & new_n15559;
  assign new_n15590 = ~new_n14949 & new_n15559;
  assign new_n15591 = ~new_n14956 & new_n15559;
  assign new_n15592 = ~new_n8448 & new_n8513;
  assign new_n15593 = ~new_n9310 & new_n15592;
  assign new_n15594 = ~new_n10088 & new_n15592;
  assign new_n15595 = ~new_n10870 & new_n15592;
  assign new_n15596 = ~new_n11648 & new_n15592;
  assign new_n15597 = ~new_n12426 & new_n15592;
  assign new_n15598 = ~new_n13204 & new_n15592;
  assign new_n15599 = ~new_n13982 & new_n15592;
  assign new_n15600 = ~new_n14760 & new_n15592;
  assign new_n15601 = ~new_n14771 & new_n15592;
  assign new_n15602 = ~new_n14781 & new_n15592;
  assign new_n15603 = ~new_n14791 & new_n15592;
  assign new_n15604 = ~new_n14801 & new_n15592;
  assign new_n15605 = ~new_n14811 & new_n15592;
  assign new_n15606 = ~new_n14821 & new_n15592;
  assign new_n15607 = ~new_n14831 & new_n15592;
  assign new_n15608 = ~new_n14841 & new_n15592;
  assign new_n15609 = ~new_n14851 & new_n15592;
  assign new_n15610 = ~new_n14858 & new_n15592;
  assign new_n15611 = ~new_n14865 & new_n15592;
  assign new_n15612 = ~new_n14872 & new_n15592;
  assign new_n15613 = ~new_n14879 & new_n15592;
  assign new_n15614 = ~new_n14886 & new_n15592;
  assign new_n15615 = ~new_n14893 & new_n15592;
  assign new_n15616 = ~new_n14900 & new_n15592;
  assign new_n15617 = ~new_n14907 & new_n15592;
  assign new_n15618 = ~new_n14914 & new_n15592;
  assign new_n15619 = ~new_n14921 & new_n15592;
  assign new_n15620 = ~new_n14928 & new_n15592;
  assign new_n15621 = ~new_n14935 & new_n15592;
  assign new_n15622 = ~new_n14942 & new_n15592;
  assign new_n15623 = ~new_n14949 & new_n15592;
  assign new_n15624 = ~new_n14956 & new_n15592;
  assign new_n15625 = ~new_n8448 & new_n14958;
  assign new_n15626 = ~new_n9310 & new_n15625;
  assign new_n15627 = ~new_n10088 & new_n15625;
  assign new_n15628 = ~new_n10870 & new_n15625;
  assign new_n15629 = ~new_n11648 & new_n15625;
  assign new_n15630 = ~new_n12426 & new_n15625;
  assign new_n15631 = ~new_n13204 & new_n15625;
  assign new_n15632 = ~new_n13982 & new_n15625;
  assign new_n15633 = ~new_n14760 & new_n15625;
  assign new_n15634 = ~new_n14771 & new_n15625;
  assign new_n15635 = ~new_n14781 & new_n15625;
  assign new_n15636 = ~new_n14791 & new_n15625;
  assign new_n15637 = ~new_n14801 & new_n15625;
  assign new_n15638 = ~new_n14811 & new_n15625;
  assign new_n15639 = ~new_n14821 & new_n15625;
  assign new_n15640 = ~new_n14831 & new_n15625;
  assign new_n15641 = ~new_n14841 & new_n15625;
  assign new_n15642 = ~new_n14851 & new_n15625;
  assign new_n15643 = ~new_n14858 & new_n15625;
  assign new_n15644 = ~new_n14865 & new_n15625;
  assign new_n15645 = ~new_n14872 & new_n15625;
  assign new_n15646 = ~new_n14879 & new_n15625;
  assign new_n15647 = ~new_n14886 & new_n15625;
  assign new_n15648 = ~new_n14893 & new_n15625;
  assign new_n15649 = ~new_n14900 & new_n15625;
  assign new_n15650 = ~new_n14907 & new_n15625;
  assign new_n15651 = ~new_n14914 & new_n15625;
  assign new_n15652 = ~new_n14921 & new_n15625;
  assign new_n15653 = ~new_n14928 & new_n15625;
  assign new_n15654 = ~new_n14935 & new_n15625;
  assign new_n15655 = ~new_n14942 & new_n15625;
  assign new_n15656 = ~new_n14949 & new_n15625;
  assign new_n15657 = ~new_n14956 & new_n15625;
  assign new_n15658 = ~new_n8448 & new_n14993;
  assign new_n15659 = ~new_n9310 & new_n15658;
  assign new_n15660 = ~new_n10088 & new_n15658;
  assign new_n15661 = ~new_n10870 & new_n15658;
  assign new_n15662 = ~new_n11648 & new_n15658;
  assign new_n15663 = ~new_n12426 & new_n15658;
  assign new_n15664 = ~new_n13204 & new_n15658;
  assign new_n15665 = ~new_n13982 & new_n15658;
  assign new_n15666 = ~new_n14760 & new_n15658;
  assign new_n15667 = ~new_n14771 & new_n15658;
  assign new_n15668 = ~new_n14781 & new_n15658;
  assign new_n15669 = ~new_n14791 & new_n15658;
  assign new_n15670 = ~new_n14801 & new_n15658;
  assign new_n15671 = ~new_n14811 & new_n15658;
  assign new_n15672 = ~new_n14821 & new_n15658;
  assign new_n15673 = ~new_n14831 & new_n15658;
  assign new_n15674 = ~new_n14841 & new_n15658;
  assign new_n15675 = ~new_n14851 & new_n15658;
  assign new_n15676 = ~new_n14858 & new_n15658;
  assign new_n15677 = ~new_n14865 & new_n15658;
  assign new_n15678 = ~new_n14872 & new_n15658;
  assign new_n15679 = ~new_n14879 & new_n15658;
  assign new_n15680 = ~new_n14886 & new_n15658;
  assign new_n15681 = ~new_n14893 & new_n15658;
  assign new_n15682 = ~new_n14900 & new_n15658;
  assign new_n15683 = ~new_n14907 & new_n15658;
  assign new_n15684 = ~new_n14914 & new_n15658;
  assign new_n15685 = ~new_n14921 & new_n15658;
  assign new_n15686 = ~new_n14928 & new_n15658;
  assign new_n15687 = ~new_n14935 & new_n15658;
  assign new_n15688 = ~new_n14942 & new_n15658;
  assign new_n15689 = ~new_n14949 & new_n15658;
  assign new_n15690 = ~new_n14956 & new_n15658;
  assign new_n15691 = new_n8447 & new_n15028;
  assign new_n15692 = ~new_n9310 & new_n15691;
  assign new_n15693 = ~new_n10088 & new_n15691;
  assign new_n15694 = ~new_n10870 & new_n15691;
  assign new_n15695 = ~new_n11648 & new_n15691;
  assign new_n15696 = ~new_n12426 & new_n15691;
  assign new_n15697 = ~new_n13204 & new_n15691;
  assign new_n15698 = ~new_n13982 & new_n15691;
  assign new_n15699 = ~new_n14760 & new_n15691;
  assign new_n15700 = ~new_n14771 & new_n15691;
  assign new_n15701 = ~new_n14781 & new_n15691;
  assign new_n15702 = ~new_n14791 & new_n15691;
  assign new_n15703 = ~new_n14801 & new_n15691;
  assign new_n15704 = ~new_n14811 & new_n15691;
  assign new_n15705 = ~new_n14821 & new_n15691;
  assign new_n15706 = ~new_n14831 & new_n15691;
  assign new_n15707 = ~new_n14841 & new_n15691;
  assign new_n15708 = ~new_n14851 & new_n15691;
  assign new_n15709 = ~new_n14858 & new_n15691;
  assign new_n15710 = ~new_n14865 & new_n15691;
  assign new_n15711 = ~new_n14872 & new_n15691;
  assign new_n15712 = ~new_n14879 & new_n15691;
  assign new_n15713 = ~new_n14886 & new_n15691;
  assign new_n15714 = ~new_n14893 & new_n15691;
  assign new_n15715 = ~new_n14900 & new_n15691;
  assign new_n15716 = ~new_n14907 & new_n15691;
  assign new_n15717 = ~new_n14914 & new_n15691;
  assign new_n15718 = ~new_n14921 & new_n15691;
  assign new_n15719 = ~new_n14928 & new_n15691;
  assign new_n15720 = ~new_n14935 & new_n15691;
  assign new_n15721 = ~new_n14942 & new_n15691;
  assign new_n15722 = ~new_n14949 & new_n15691;
  assign new_n15723 = ~new_n14956 & new_n15691;
  assign new_n15724 = new_n8447 & new_n8514;
  assign new_n15725 = ~new_n9310 & new_n15724;
  assign new_n15726 = ~new_n10088 & new_n15724;
  assign new_n15727 = ~new_n10870 & new_n15724;
  assign new_n15728 = ~new_n11648 & new_n15724;
  assign new_n15729 = ~new_n12426 & new_n15724;
  assign new_n15730 = ~new_n13204 & new_n15724;
  assign new_n15731 = ~new_n13982 & new_n15724;
  assign new_n15732 = ~new_n14760 & new_n15724;
  assign new_n15733 = ~new_n14771 & new_n15724;
  assign new_n15734 = ~new_n14781 & new_n15724;
  assign new_n15735 = ~new_n14791 & new_n15724;
  assign new_n15736 = ~new_n14801 & new_n15724;
  assign new_n15737 = ~new_n14811 & new_n15724;
  assign new_n15738 = ~new_n14821 & new_n15724;
  assign new_n15739 = ~new_n14831 & new_n15724;
  assign new_n15740 = ~new_n14841 & new_n15724;
  assign new_n15741 = ~new_n14851 & new_n15724;
  assign new_n15742 = ~new_n14858 & new_n15724;
  assign new_n15743 = ~new_n14865 & new_n15724;
  assign new_n15744 = ~new_n14872 & new_n15724;
  assign new_n15745 = ~new_n14879 & new_n15724;
  assign new_n15746 = ~new_n14886 & new_n15724;
  assign new_n15747 = ~new_n14893 & new_n15724;
  assign new_n15748 = ~new_n14900 & new_n15724;
  assign new_n15749 = ~new_n14907 & new_n15724;
  assign new_n15750 = ~new_n14914 & new_n15724;
  assign new_n15751 = ~new_n14921 & new_n15724;
  assign new_n15752 = ~new_n14928 & new_n15724;
  assign new_n15753 = ~new_n14935 & new_n15724;
  assign new_n15754 = ~new_n14942 & new_n15724;
  assign new_n15755 = ~new_n14949 & new_n15724;
  assign new_n15756 = ~new_n14956 & new_n15724;
  assign new_n15757 = new_n8447 & new_n14959;
  assign new_n15758 = ~new_n9310 & new_n15757;
  assign new_n15759 = ~new_n10088 & new_n15757;
  assign new_n15760 = ~new_n10870 & new_n15757;
  assign new_n15761 = ~new_n11648 & new_n15757;
  assign new_n15762 = ~new_n12426 & new_n15757;
  assign new_n15763 = ~new_n13204 & new_n15757;
  assign new_n15764 = ~new_n13982 & new_n15757;
  assign new_n15765 = ~new_n14760 & new_n15757;
  assign new_n15766 = ~new_n14771 & new_n15757;
  assign new_n15767 = ~new_n14781 & new_n15757;
  assign new_n15768 = ~new_n14791 & new_n15757;
  assign new_n15769 = ~new_n14801 & new_n15757;
  assign new_n15770 = ~new_n14811 & new_n15757;
  assign new_n15771 = ~new_n14821 & new_n15757;
  assign new_n15772 = ~new_n14831 & new_n15757;
  assign new_n15773 = ~new_n14841 & new_n15757;
  assign new_n15774 = ~new_n14851 & new_n15757;
  assign new_n15775 = ~new_n14858 & new_n15757;
  assign new_n15776 = ~new_n14865 & new_n15757;
  assign new_n15777 = ~new_n14872 & new_n15757;
  assign new_n15778 = ~new_n14879 & new_n15757;
  assign new_n15779 = ~new_n14886 & new_n15757;
  assign new_n15780 = ~new_n14893 & new_n15757;
  assign new_n15781 = ~new_n14900 & new_n15757;
  assign new_n15782 = ~new_n14907 & new_n15757;
  assign new_n15783 = ~new_n14914 & new_n15757;
  assign new_n15784 = ~new_n14921 & new_n15757;
  assign new_n15785 = ~new_n14928 & new_n15757;
  assign new_n15786 = ~new_n14935 & new_n15757;
  assign new_n15787 = ~new_n14942 & new_n15757;
  assign new_n15788 = ~new_n14949 & new_n15757;
  assign new_n15789 = ~new_n14956 & new_n15757;
  assign new_n15790 = ~new_n14994 & new_n8447;
  assign new_n15791 = ~new_n9310 & new_n15790;
  assign new_n15792 = ~new_n10088 & new_n15790;
  assign new_n15793 = ~new_n10870 & new_n15790;
  assign new_n15794 = ~new_n11648 & new_n15790;
  assign new_n15795 = ~new_n12426 & new_n15790;
  assign new_n15796 = ~new_n13204 & new_n15790;
  assign new_n15797 = ~new_n13982 & new_n15790;
  assign new_n15798 = ~new_n14760 & new_n15790;
  assign new_n15799 = ~new_n14771 & new_n15790;
  assign new_n15800 = ~new_n14781 & new_n15790;
  assign new_n15801 = ~new_n14791 & new_n15790;
  assign new_n15802 = ~new_n14801 & new_n15790;
  assign new_n15803 = ~new_n14811 & new_n15790;
  assign new_n15804 = ~new_n14821 & new_n15790;
  assign new_n15805 = ~new_n14831 & new_n15790;
  assign new_n15806 = ~new_n14841 & new_n15790;
  assign new_n15807 = ~new_n14851 & new_n15790;
  assign new_n15808 = ~new_n14858 & new_n15790;
  assign new_n15809 = ~new_n14865 & new_n15790;
  assign new_n15810 = ~new_n14872 & new_n15790;
  assign new_n15811 = ~new_n14879 & new_n15790;
  assign new_n15812 = ~new_n14886 & new_n15790;
  assign new_n15813 = ~new_n14893 & new_n15790;
  assign new_n15814 = ~new_n14900 & new_n15790;
  assign new_n15815 = ~new_n14907 & new_n15790;
  assign new_n15816 = ~new_n14914 & new_n15790;
  assign new_n15817 = ~new_n14921 & new_n15790;
  assign new_n15818 = ~new_n14928 & new_n15790;
  assign new_n15819 = ~new_n14935 & new_n15790;
  assign new_n15820 = ~new_n14942 & new_n15790;
  assign new_n15821 = ~new_n14949 & new_n15790;
  assign new_n15822 = ~new_n14956 & new_n15790;
  assign new_n15823 = new_n8447 & new_n15029;
  assign new_n15824 = ~new_n9310 & new_n15823;
  assign new_n15825 = ~new_n10088 & new_n15823;
  assign new_n15826 = ~new_n10870 & new_n15823;
  assign new_n15827 = ~new_n11648 & new_n15823;
  assign new_n15828 = ~new_n12426 & new_n15823;
  assign new_n15829 = ~new_n13204 & new_n15823;
  assign new_n15830 = ~new_n13982 & new_n15823;
  assign new_n15831 = ~new_n14760 & new_n15823;
  assign new_n15832 = ~new_n14771 & new_n15823;
  assign new_n15833 = ~new_n14781 & new_n15823;
  assign new_n15834 = ~new_n14791 & new_n15823;
  assign new_n15835 = ~new_n14801 & new_n15823;
  assign new_n15836 = ~new_n14811 & new_n15823;
  assign new_n15837 = ~new_n14821 & new_n15823;
  assign new_n15838 = ~new_n14831 & new_n15823;
  assign new_n15839 = ~new_n14841 & new_n15823;
  assign new_n15840 = ~new_n14851 & new_n15823;
  assign new_n15841 = ~new_n14858 & new_n15823;
  assign new_n15842 = ~new_n14865 & new_n15823;
  assign new_n15843 = ~new_n14872 & new_n15823;
  assign new_n15844 = ~new_n14879 & new_n15823;
  assign new_n15845 = ~new_n14886 & new_n15823;
  assign new_n15846 = ~new_n14893 & new_n15823;
  assign new_n15847 = ~new_n14900 & new_n15823;
  assign new_n15848 = ~new_n14907 & new_n15823;
  assign new_n15849 = ~new_n14914 & new_n15823;
  assign new_n15850 = ~new_n14921 & new_n15823;
  assign new_n15851 = ~new_n14928 & new_n15823;
  assign new_n15852 = ~new_n14935 & new_n15823;
  assign new_n15853 = ~new_n14942 & new_n15823;
  assign new_n15854 = ~new_n14949 & new_n15823;
  assign new_n15855 = ~new_n14956 & new_n15823;
  assign new_n15856 = new_n8447 & new_n8513;
  assign new_n15857 = ~new_n9310 & new_n15856;
  assign new_n15858 = ~new_n10088 & new_n15856;
  assign new_n15859 = ~new_n10870 & new_n15856;
  assign new_n15860 = ~new_n11648 & new_n15856;
  assign new_n15861 = ~new_n12426 & new_n15856;
  assign new_n15862 = ~new_n13204 & new_n15856;
  assign new_n15863 = ~new_n13982 & new_n15856;
  assign new_n15864 = ~new_n14760 & new_n15856;
  assign new_n15865 = ~new_n14771 & new_n15856;
  assign new_n15866 = ~new_n14781 & new_n15856;
  assign new_n15867 = ~new_n14791 & new_n15856;
  assign new_n15868 = ~new_n14801 & new_n15856;
  assign new_n15869 = ~new_n14811 & new_n15856;
  assign new_n15870 = ~new_n14821 & new_n15856;
  assign new_n15871 = ~new_n14831 & new_n15856;
  assign new_n15872 = ~new_n14841 & new_n15856;
  assign new_n15873 = ~new_n14851 & new_n15856;
  assign new_n15874 = ~new_n14858 & new_n15856;
  assign new_n15875 = ~new_n14865 & new_n15856;
  assign new_n15876 = ~new_n14872 & new_n15856;
  assign new_n15877 = ~new_n14879 & new_n15856;
  assign new_n15878 = ~new_n14886 & new_n15856;
  assign new_n15879 = ~new_n14893 & new_n15856;
  assign new_n15880 = ~new_n14900 & new_n15856;
  assign new_n15881 = ~new_n14907 & new_n15856;
  assign new_n15882 = ~new_n14914 & new_n15856;
  assign new_n15883 = ~new_n14921 & new_n15856;
  assign new_n15884 = ~new_n14928 & new_n15856;
  assign new_n15885 = ~new_n14935 & new_n15856;
  assign new_n15886 = ~new_n14942 & new_n15856;
  assign new_n15887 = ~new_n14949 & new_n15856;
  assign new_n15888 = ~new_n14956 & new_n15856;
  assign new_n15889 = new_n8447 & new_n14958;
  assign new_n15890 = ~new_n9310 & new_n15889;
  assign new_n15891 = ~new_n10088 & new_n15889;
  assign new_n15892 = ~new_n10870 & new_n15889;
  assign new_n15893 = ~new_n11648 & new_n15889;
  assign new_n15894 = ~new_n12426 & new_n15889;
  assign new_n15895 = ~new_n13204 & new_n15889;
  assign new_n15896 = ~new_n13982 & new_n15889;
  assign new_n15897 = ~new_n14760 & new_n15889;
  assign new_n15898 = ~new_n14771 & new_n15889;
  assign new_n15899 = ~new_n14781 & new_n15889;
  assign new_n15900 = ~new_n14791 & new_n15889;
  assign new_n15901 = ~new_n14801 & new_n15889;
  assign new_n15902 = ~new_n14811 & new_n15889;
  assign new_n15903 = ~new_n14821 & new_n15889;
  assign new_n15904 = ~new_n14831 & new_n15889;
  assign new_n15905 = ~new_n14841 & new_n15889;
  assign new_n15906 = ~new_n14851 & new_n15889;
  assign new_n15907 = ~new_n14858 & new_n15889;
  assign new_n15908 = ~new_n14865 & new_n15889;
  assign new_n15909 = ~new_n14872 & new_n15889;
  assign new_n15910 = ~new_n14879 & new_n15889;
  assign new_n15911 = ~new_n14886 & new_n15889;
  assign new_n15912 = ~new_n14893 & new_n15889;
  assign new_n15913 = ~new_n14900 & new_n15889;
  assign new_n15914 = ~new_n14907 & new_n15889;
  assign new_n15915 = ~new_n14914 & new_n15889;
  assign new_n15916 = ~new_n14921 & new_n15889;
  assign new_n15917 = ~new_n14928 & new_n15889;
  assign new_n15918 = ~new_n14935 & new_n15889;
  assign new_n15919 = ~new_n14942 & new_n15889;
  assign new_n15920 = ~new_n14949 & new_n15889;
  assign new_n15921 = ~new_n14956 & new_n15889;
  assign new_n15922 = new_n8447 & new_n14993;
  assign new_n15923 = ~new_n9310 & new_n15922;
  assign new_n15924 = ~new_n10088 & new_n15922;
  assign new_n15925 = ~new_n10870 & new_n15922;
  assign new_n15926 = ~new_n11648 & new_n15922;
  assign new_n15927 = ~new_n12426 & new_n15922;
  assign new_n15928 = ~new_n13204 & new_n15922;
  assign new_n15929 = ~new_n13982 & new_n15922;
  assign new_n15930 = ~new_n14760 & new_n15922;
  assign new_n15931 = ~new_n14771 & new_n15922;
  assign new_n15932 = ~new_n14781 & new_n15922;
  assign new_n15933 = ~new_n14791 & new_n15922;
  assign new_n15934 = ~new_n14801 & new_n15922;
  assign new_n15935 = ~new_n14811 & new_n15922;
  assign new_n15936 = ~new_n14821 & new_n15922;
  assign new_n15937 = ~new_n14831 & new_n15922;
  assign new_n15938 = ~new_n14841 & new_n15922;
  assign new_n15939 = ~new_n14851 & new_n15922;
  assign new_n15940 = ~new_n14858 & new_n15922;
  assign new_n15941 = ~new_n14865 & new_n15922;
  assign new_n15942 = ~new_n14872 & new_n15922;
  assign new_n15943 = ~new_n14879 & new_n15922;
  assign new_n15944 = ~new_n14886 & new_n15922;
  assign new_n15945 = ~new_n14893 & new_n15922;
  assign new_n15946 = ~new_n14900 & new_n15922;
  assign new_n15947 = ~new_n14907 & new_n15922;
  assign new_n15948 = ~new_n14914 & new_n15922;
  assign new_n15949 = ~new_n14921 & new_n15922;
  assign new_n15950 = ~new_n14928 & new_n15922;
  assign new_n15951 = ~new_n14935 & new_n15922;
  assign new_n15952 = ~new_n14942 & new_n15922;
  assign new_n15953 = ~new_n14949 & new_n15922;
  assign new_n15954 = ~new_n14956 & new_n15922;
  assign po0 = n2049;
  assign po1 = n2050;
  assign po2 = n2051;
  assign po3 = n2052;
  assign po4 = n2053;
  assign po5 = n2054;
  assign po6 = n2055;
  assign po7 = n2056;
  assign po8 = n2057;
  assign po9 = n2058;
  assign po10 = n2059;
  assign po11 = n2060;
  assign po12 = n2061;
  assign po13 = n2062;
  assign po14 = n2063;
  assign po15 = n2064;
  assign po16 = n2065;
  assign po17 = n2066;
  assign po18 = n2067;
  assign po19 = n2068;
  assign po20 = n2069;
  assign po21 = n2070;
  assign po22 = n2071;
  assign po23 = n2072;
  assign po24 = n2073;
  assign po25 = n2074;
  assign po26 = n2075;
  assign po27 = n2076;
  assign po28 = n2077;
  assign po29 = n2078;
  assign po30 = n2079;
  assign po31 = n2080;
  assign po32 = n2081;
  assign po33 = n2082;
  assign po34 = n2083;
  assign po35 = n2084;
  assign po36 = n2085;
  assign po37 = n2086;
  assign po38 = n2087;
  assign po39 = n2088;
  assign po40 = n2089;
  assign po41 = n2090;
  assign po42 = n2091;
  assign po43 = n2092;
  assign po44 = n2093;
  assign po45 = n2094;
  assign po46 = n2095;
  assign po47 = n2096;
  assign po48 = n2097;
  assign po49 = n2098;
  assign po50 = n2099;
  assign po51 = n2100;
  assign po52 = n2101;
  assign po53 = n2102;
  assign po54 = n2103;
  assign po55 = n2104;
  assign po56 = n2105;
  assign po57 = n2106;
  assign po58 = n2107;
  assign po59 = n2108;
  assign po60 = n2109;
  assign po61 = n2110;
  assign po62 = n2111;
  assign po63 = n2112;
  assign po64 = n2113;
  assign po65 = n2114;
  assign po66 = n2115;
  assign po67 = n2116;
  assign po68 = n2117;
  assign po69 = n2118;
  assign po70 = n2119;
  assign po71 = n2120;
  assign po72 = n2121;
  assign po73 = n2122;
  assign po74 = n2123;
  assign po75 = n2124;
  assign po76 = n2125;
  assign po77 = n2126;
  assign po78 = n2127;
  assign po79 = n2128;
  assign po80 = n2129;
  assign po81 = n2130;
  assign po82 = n2131;
  assign po83 = n2132;
  assign po84 = n2133;
  assign po85 = n2134;
  assign po86 = n2135;
  assign po87 = n2136;
  assign po88 = n2137;
  assign po89 = n2138;
  assign po90 = n2139;
  assign po91 = n2140;
  assign po92 = n2141;
  assign po93 = n2142;
  assign po94 = n2143;
  assign po95 = n2144;
  assign po96 = n2145;
  assign po97 = n2146;
  assign po98 = n2147;
  assign po99 = n2148;
  assign po100 = n2149;
  assign po101 = n2150;
  assign po102 = n2151;
  assign po103 = n2152;
  assign po104 = n2153;
  assign po105 = n2154;
  assign po106 = n2155;
  assign po107 = n2156;
  assign po108 = n2157;
  assign po109 = n2158;
  assign po110 = n2159;
  assign po111 = n2160;
  assign po112 = n2161;
  assign po113 = n2162;
  assign po114 = n2163;
  assign po115 = n2164;
  assign po116 = n2165;
  assign po117 = n2166;
  assign po118 = n2167;
  assign po119 = n2168;
  assign po120 = n2169;
  assign po121 = n2170;
  assign po122 = n2171;
  assign po123 = n2172;
  assign po124 = n2173;
  assign po125 = n2174;
  assign po126 = n2175;
  assign po127 = n2176;
  assign po128 = n2177;
  assign po129 = n2178;
  assign po130 = n2179;
  assign po131 = n2180;
  assign po132 = n2181;
  assign po133 = n2182;
  assign po134 = n2183;
  assign po135 = n2184;
  assign po136 = n2185;
  assign po137 = n2186;
  assign po138 = n2187;
  assign po139 = n2188;
  assign po140 = n2189;
  assign po141 = n2190;
  assign po142 = n2191;
  assign po143 = n2192;
  assign po144 = n2193;
  assign po145 = n2194;
  assign po146 = n2195;
  assign po147 = n2196;
  assign po148 = n2197;
  assign po149 = n2198;
  assign po150 = n2199;
  assign po151 = n2200;
  assign po152 = n2201;
  assign po153 = n2202;
  assign po154 = n2203;
  assign po155 = n2204;
  assign po156 = n2205;
  assign po157 = n2206;
  assign po158 = n2207;
  assign po159 = n2208;
  assign po160 = n2209;
  assign po161 = n2210;
  assign po162 = n2211;
  assign po163 = n2212;
  assign po164 = n2213;
  assign po165 = n2214;
  assign po166 = n2215;
  assign po167 = n2216;
  assign po168 = n2217;
  assign po169 = n2218;
  assign po170 = n2219;
  assign po171 = n2220;
  assign po172 = n2221;
  assign po173 = n2222;
  assign po174 = n2223;
  assign po175 = n2224;
  assign po176 = n2225;
  assign po177 = n2226;
  assign po178 = n2227;
  assign po179 = n2228;
  assign po180 = n2229;
  assign po181 = n2230;
  assign po182 = n2231;
  assign po183 = n2232;
  assign po184 = n2233;
  assign po185 = n2234;
  assign po186 = n2235;
  assign po187 = n2236;
  assign po188 = n2237;
  assign po189 = n2238;
  assign po190 = n2239;
  assign po191 = n2240;
  assign po192 = n2241;
  assign po193 = n2242;
  assign po194 = n2243;
  assign po195 = n2244;
  assign po196 = n2245;
  assign po197 = n2246;
  assign po198 = n2247;
  assign po199 = n2248;
  assign po200 = n2249;
  assign po201 = n2250;
  assign po202 = n2251;
  assign po203 = n2252;
  assign po204 = n2253;
  assign po205 = n2254;
  assign po206 = n2255;
  assign po207 = n2256;
  assign po208 = n2257;
  assign po209 = n2258;
  assign po210 = n2259;
  assign po211 = n2260;
  assign po212 = n2261;
  assign po213 = n2262;
  assign po214 = n2263;
  assign po215 = n2264;
  assign po216 = n2265;
  assign po217 = n2266;
  assign po218 = n2267;
  assign po219 = n2268;
  assign po220 = n2269;
  assign po221 = n2270;
  assign po222 = n2271;
  assign po223 = n2272;
  assign po224 = n2273;
  assign po225 = n2274;
  assign po226 = n2275;
  assign po227 = n2276;
  assign po228 = n2277;
  assign po229 = n2278;
  assign po230 = n2279;
  assign po231 = n2280;
  assign po232 = n2281;
  assign po233 = n2282;
  assign po234 = n2283;
  assign po235 = n2284;
  assign po236 = n2285;
  assign po237 = n2286;
  assign po238 = n2287;
  assign po239 = n2288;
  assign po240 = n2289;
  assign po241 = n2290;
  assign po242 = n2291;
  assign po243 = n2292;
  assign po244 = n2293;
  assign po245 = n2294;
  assign po246 = n2295;
  assign po247 = n2296;
  assign po248 = n2297;
  assign po249 = n2298;
  assign po250 = n2299;
  assign po251 = n2300;
  assign po252 = n2301;
  assign po253 = n2302;
  assign po254 = n2303;
  assign po255 = n2304;
  assign po256 = n2305;
  assign po257 = n2306;
  assign po258 = n2307;
  assign po259 = n2308;
  assign po260 = n2309;
  assign po261 = n2310;
  assign po262 = n2311;
  assign po263 = n2312;
  assign po264 = n2313;
  assign po265 = n2314;
  assign po266 = n2315;
  assign po267 = n2316;
  assign po268 = n2317;
  assign po269 = n2318;
  assign po270 = n2319;
  assign po271 = n2320;
  assign po272 = n2321;
  assign po273 = n2322;
  assign po274 = n2323;
  assign po275 = n2324;
  assign po276 = n2325;
  assign po277 = n2326;
  assign po278 = n2327;
  assign po279 = n2328;
  assign po280 = n2329;
  assign po281 = n2330;
  assign po282 = n2331;
  assign po283 = n2332;
  assign po284 = n2333;
  assign po285 = n2334;
  assign po286 = n2335;
  assign po287 = n2336;
  assign po288 = n2337;
  assign po289 = n2338;
  assign po290 = n2339;
  assign po291 = n2340;
  assign po292 = n2341;
  assign po293 = n2342;
  assign po294 = n2343;
  assign po295 = n2344;
  assign po296 = n2345;
  assign po297 = n2346;
  assign po298 = n2347;
  assign po299 = n2348;
  assign po300 = n2349;
  assign po301 = n2350;
  assign po302 = n2351;
  assign po303 = n2352;
  assign po304 = n2353;
  assign po305 = n2354;
  assign po306 = n2355;
  assign po307 = n2356;
  assign po308 = n2357;
  assign po309 = n2358;
  assign po310 = n2359;
  assign po311 = n2360;
  assign po312 = n2361;
  assign po313 = n2362;
  assign po314 = n2363;
  assign po315 = n2364;
  assign po316 = n2365;
  assign po317 = n2366;
  assign po318 = n2367;
  assign po319 = n2368;
  assign po320 = n2369;
  assign po321 = n2370;
  assign po322 = n2371;
  assign po323 = n2372;
  assign po324 = n2373;
  assign po325 = n2374;
  assign po326 = n2375;
  assign po327 = n2376;
  assign po328 = n2377;
  assign po329 = n2378;
  assign po330 = n2379;
  assign po331 = n2380;
  assign po332 = n2381;
  assign po333 = n2382;
  assign po334 = n2383;
  assign po335 = n2384;
  assign po336 = n2385;
  assign po337 = n2386;
  assign po338 = n2387;
  assign po339 = n2388;
  assign po340 = n2389;
  assign po341 = n2390;
  assign po342 = n2391;
  assign po343 = n2392;
  assign po344 = n2393;
  assign po345 = n2394;
  assign po346 = n2395;
  assign po347 = n2396;
  assign po348 = n2397;
  assign po349 = n2398;
  assign po350 = n2399;
  assign po351 = n2400;
  assign po352 = n2401;
  assign po353 = n2402;
  assign po354 = n2403;
  assign po355 = n2404;
  assign po356 = n2405;
  assign po357 = n2406;
  assign po358 = n2407;
  assign po359 = n2408;
  assign po360 = n2409;
  assign po361 = n2410;
  assign po362 = n2411;
  assign po363 = n2412;
  assign po364 = n2413;
  assign po365 = n2414;
  assign po366 = n2415;
  assign po367 = n2416;
  assign po368 = n2417;
  assign po369 = n2418;
  assign po370 = n2419;
  assign po371 = n2420;
  assign po372 = n2421;
  assign po373 = n2422;
  assign po374 = n2423;
  assign po375 = n2424;
  assign po376 = n2425;
  assign po377 = n2426;
  assign po378 = n2427;
  assign po379 = n2428;
  assign po380 = n2429;
  assign po381 = n2430;
  assign po382 = n2431;
  assign po383 = n2432;
  assign po384 = n2433;
  assign po385 = n2434;
  assign po386 = n2435;
  assign po387 = n2436;
  assign po388 = n2437;
  assign po389 = n2438;
  assign po390 = n2439;
  assign po391 = n2440;
  assign po392 = n2441;
  assign po393 = n2442;
  assign po394 = n2443;
  assign po395 = n2444;
  assign po396 = n2445;
  assign po397 = n2446;
  assign po398 = n2447;
  assign po399 = n2448;
  assign po400 = n2449;
  assign po401 = n2450;
  assign po402 = n2451;
  assign po403 = n2452;
  assign po404 = n2453;
  assign po405 = n2454;
  assign po406 = n2455;
  assign po407 = n2456;
  assign po408 = n2457;
  assign po409 = n2458;
  assign po410 = n2459;
  assign po411 = n2460;
  assign po412 = n2461;
  assign po413 = n2462;
  assign po414 = n2463;
  assign po415 = n2464;
  assign po416 = n2465;
  assign po417 = n2466;
  assign po418 = n2467;
  assign po419 = n2468;
  assign po420 = n2469;
  assign po421 = n2470;
  assign po422 = n2471;
  assign po423 = n2472;
  assign po424 = n2473;
  assign po425 = n2474;
  assign po426 = n2475;
  assign po427 = n2476;
  assign po428 = n2477;
  assign po429 = n2478;
  assign po430 = n2479;
  assign po431 = n2480;
  assign po432 = n2481;
  assign po433 = n2482;
  assign po434 = n2483;
  assign po435 = n2484;
  assign po436 = n2485;
  assign po437 = n2486;
  assign po438 = n2487;
  assign po439 = n2488;
  assign po440 = n2489;
  assign po441 = n2490;
  assign po442 = n2491;
  assign po443 = n2492;
  assign po444 = n2493;
  assign po445 = n2494;
  assign po446 = n2495;
  assign po447 = n2496;
  assign po448 = n2497;
  assign po449 = n2498;
  assign po450 = n2499;
  assign po451 = n2500;
  assign po452 = n2501;
  assign po453 = n2502;
  assign po454 = n2503;
  assign po455 = n2504;
  assign po456 = n2505;
  assign po457 = n2506;
  assign po458 = n2507;
  assign po459 = n2508;
  assign po460 = n2509;
  assign po461 = n2510;
  assign po462 = n2511;
  assign po463 = n2512;
  assign po464 = n2513;
  assign po465 = n2514;
  assign po466 = n2515;
  assign po467 = n2516;
  assign po468 = n2517;
  assign po469 = n2518;
  assign po470 = n2519;
  assign po471 = n2520;
  assign po472 = n2521;
  assign po473 = n2522;
  assign po474 = n2523;
  assign po475 = n2524;
  assign po476 = n2525;
  assign po477 = n2526;
  assign po478 = n2527;
  assign po479 = n2528;
  assign po480 = n2529;
  assign po481 = n2530;
  assign po482 = n2531;
  assign po483 = n2532;
  assign po484 = n2533;
  assign po485 = n2534;
  assign po486 = n2535;
  assign po487 = n2536;
  assign po488 = n2537;
  assign po489 = n2538;
  assign po490 = n2539;
  assign po491 = n2540;
  assign po492 = n2541;
  assign po493 = n2542;
  assign po494 = n2543;
  assign po495 = n2544;
  assign po496 = n2545;
  assign po497 = n2546;
  assign po498 = n2547;
  assign po499 = n2548;
  assign po500 = n2549;
  assign po501 = n2550;
  assign po502 = n2551;
  assign po503 = n2552;
  assign po504 = n2553;
  assign po505 = n2554;
  assign po506 = n2555;
  assign po507 = n2556;
  assign po508 = n2557;
  assign po509 = n2558;
  assign po510 = n2559;
  assign po511 = n2560;
  assign po512 = n2561;
  assign po513 = n2562;
  assign po514 = n2563;
  assign po515 = n2564;
  assign po516 = n2565;
  assign po517 = n2566;
  assign po518 = n2567;
  assign po519 = n2568;
  assign po520 = n2569;
  assign po521 = n2570;
  assign po522 = n2571;
  assign po523 = n2572;
  assign po524 = n2573;
  assign po525 = n2574;
  assign po526 = n2575;
  assign po527 = n2576;
  assign po528 = n2577;
  assign po529 = n2578;
  assign po530 = n2579;
  assign po531 = n2580;
  assign po532 = n2581;
  assign po533 = n2582;
  assign po534 = n2583;
  assign po535 = n2584;
  assign po536 = n2585;
  assign po537 = n2586;
  assign po538 = n2587;
  assign po539 = n2588;
  assign po540 = n2589;
  assign po541 = n2590;
  assign po542 = n2591;
  assign po543 = n2592;
  assign po544 = n2593;
  assign po545 = n2594;
  assign po546 = n2595;
  assign po547 = n2596;
  assign po548 = n2597;
  assign po549 = n2598;
  assign po550 = n2599;
  assign po551 = n2600;
  assign po552 = n2601;
  assign po553 = n2602;
  assign po554 = n2603;
  assign po555 = n2604;
  assign po556 = n2605;
  assign po557 = n2606;
  assign po558 = n2607;
  assign po559 = n2608;
  assign po560 = n2609;
  assign po561 = n2610;
  assign po562 = n2611;
  assign po563 = n2612;
  assign po564 = n2613;
  assign po565 = n2614;
  assign po566 = n2615;
  assign po567 = n2616;
  assign po568 = n2617;
  assign po569 = n2618;
  assign po570 = n2619;
  assign po571 = n2620;
  assign po572 = n2621;
  assign po573 = n2622;
  assign po574 = n2623;
  assign po575 = n2624;
  assign po576 = n2625;
  assign po577 = n2626;
  assign po578 = n2627;
  assign po579 = n2628;
  assign po580 = n2629;
  assign po581 = n2630;
  assign po582 = n2631;
  assign po583 = n2632;
  assign po584 = n2633;
  assign po585 = n2634;
  assign po586 = n2635;
  assign po587 = n2636;
  assign po588 = n2637;
  assign po589 = n2638;
  assign po590 = n2639;
  assign po591 = n2640;
  assign po592 = n2641;
  assign po593 = n2642;
  assign po594 = n2643;
  assign po595 = n2644;
  assign po596 = n2645;
  assign po597 = n2646;
  assign po598 = n2647;
  assign po599 = n2648;
  assign po600 = n2649;
  assign po601 = n2650;
  assign po602 = n2651;
  assign po603 = n2652;
  assign po604 = n2653;
  assign po605 = n2654;
  assign po606 = n2655;
  assign po607 = n2656;
  assign po608 = n2657;
  assign po609 = n2658;
  assign po610 = n2659;
  assign po611 = n2660;
  assign po612 = n2661;
  assign po613 = n2662;
  assign po614 = n2663;
  assign po615 = n2664;
  assign po616 = n2665;
  assign po617 = n2666;
  assign po618 = n2667;
  assign po619 = n2668;
  assign po620 = n2669;
  assign po621 = n2670;
  assign po622 = n2671;
  assign po623 = n2672;
  assign po624 = n2673;
  assign po625 = n2674;
  assign po626 = n2675;
  assign po627 = n2676;
  assign po628 = n2677;
  assign po629 = n2678;
  assign po630 = n2679;
  assign po631 = n2680;
  assign po632 = n2681;
  assign po633 = n2682;
  assign po634 = n2683;
  assign po635 = n2684;
  assign po636 = n2685;
  assign po637 = n2686;
  assign po638 = n2687;
  assign po639 = n2688;
  assign po640 = n2689;
  assign po641 = n2690;
  assign po642 = n2691;
  assign po643 = n2692;
  assign po644 = n2693;
  assign po645 = n2694;
  assign po646 = n2695;
  assign po647 = n2696;
  assign po648 = n2697;
  assign po649 = n2698;
  assign po650 = n2699;
  assign po651 = n2700;
  assign po652 = n2701;
  assign po653 = n2702;
  assign po654 = n2703;
  assign po655 = n2704;
  assign po656 = n2705;
  assign po657 = n2706;
  assign po658 = n2707;
  assign po659 = n2708;
  assign po660 = n2709;
  assign po661 = n2710;
  assign po662 = n2711;
  assign po663 = n2712;
  assign po664 = n2713;
  assign po665 = n2714;
  assign po666 = n2715;
  assign po667 = n2716;
  assign po668 = n2717;
  assign po669 = n2718;
  assign po670 = n2719;
  assign po671 = n2720;
  assign po672 = n2721;
  assign po673 = n2722;
  assign po674 = n2723;
  assign po675 = n2724;
  assign po676 = n2725;
  assign po677 = n2726;
  assign po678 = n2727;
  assign po679 = n2728;
  assign po680 = n2729;
  assign po681 = n2730;
  assign po682 = n2731;
  assign po683 = n2732;
  assign po684 = n2733;
  assign po685 = n2734;
  assign po686 = n2735;
  assign po687 = n2736;
  assign po688 = n2737;
  assign po689 = n2738;
  assign po690 = n2739;
  assign po691 = n2740;
  assign po692 = n2741;
  assign po693 = n2742;
  assign po694 = n2743;
  assign po695 = n2744;
  assign po696 = n2745;
  assign po697 = n2746;
  assign po698 = n2747;
  assign po699 = n2748;
  assign po700 = n2749;
  assign po701 = n2750;
  assign po702 = n2751;
  assign po703 = n2752;
  assign po704 = n2753;
  assign po705 = n2754;
  assign po706 = n2755;
  assign po707 = n2756;
  assign po708 = n2757;
  assign po709 = n2758;
  assign po710 = n2759;
  assign po711 = n2760;
  assign po712 = n2761;
  assign po713 = n2762;
  assign po714 = n2763;
  assign po715 = n2764;
  assign po716 = n2765;
  assign po717 = n2766;
  assign po718 = n2767;
  assign po719 = n2768;
  assign po720 = n2769;
  assign po721 = n2770;
  assign po722 = n2771;
  assign po723 = n2772;
  assign po724 = n2773;
  assign po725 = n2774;
  assign po726 = n2775;
  assign po727 = n2776;
  assign po728 = n2777;
  assign po729 = n2778;
  assign po730 = n2779;
  assign po731 = n2780;
  assign po732 = n2781;
  assign po733 = n2782;
  assign po734 = n2783;
  assign po735 = n2784;
  assign po736 = n2785;
  assign po737 = n2786;
  assign po738 = n2787;
  assign po739 = n2788;
  assign po740 = n2789;
  assign po741 = n2790;
  assign po742 = n2791;
  assign po743 = n2792;
  assign po744 = n2793;
  assign po745 = n2794;
  assign po746 = n2795;
  assign po747 = n2796;
  assign po748 = n2797;
  assign po749 = n2798;
  assign po750 = n2799;
  assign po751 = n2800;
  assign po752 = n2801;
  assign po753 = n2802;
  assign po754 = n2803;
  assign po755 = n2804;
  assign po756 = n2805;
  assign po757 = n2806;
  assign po758 = n2807;
  assign po759 = n2808;
  assign po760 = n2809;
  assign po761 = n2810;
  assign po762 = n2811;
  assign po763 = n2812;
  assign po764 = n2813;
  assign po765 = n2814;
  assign po766 = n2815;
  assign po767 = n2816;
  assign po768 = n2817;
  assign po769 = n2818;
  assign po770 = n2819;
  assign po771 = n2820;
  assign po772 = n2821;
  assign po773 = n2822;
  assign po774 = n2823;
  assign po775 = n2824;
  assign po776 = n2825;
  assign po777 = n2826;
  assign po778 = n2827;
  assign po779 = n2828;
  assign po780 = n2829;
  assign po781 = n2830;
  assign po782 = n2831;
  assign po783 = n2832;
  assign po784 = n2833;
  assign po785 = n2834;
  assign po786 = n2835;
  assign po787 = n2836;
  assign po788 = n2837;
  assign po789 = n2838;
  assign po790 = n2839;
  assign po791 = n2840;
  assign po792 = n2841;
  assign po793 = n2842;
  assign po794 = n2843;
  assign po795 = n2844;
  assign po796 = n2845;
  assign po797 = n2846;
  assign po798 = n2847;
  assign po799 = n2848;
  assign po800 = n2849;
  assign po801 = n2850;
  assign po802 = n2851;
  assign po803 = n2852;
  assign po804 = n2853;
  assign po805 = n2854;
  assign po806 = n2855;
  assign po807 = n2856;
  assign po808 = n2857;
  assign po809 = n2858;
  assign po810 = n2859;
  assign po811 = n2860;
  assign po812 = n2861;
  assign po813 = n2862;
  assign po814 = n2863;
  assign po815 = n2864;
  assign po816 = n2865;
  assign po817 = n2866;
  assign po818 = n2867;
  assign po819 = n2868;
  assign po820 = n2869;
  assign po821 = n2870;
  assign po822 = n2871;
  assign po823 = n2872;
  assign po824 = n2873;
  assign po825 = n2874;
  assign po826 = n2875;
  assign po827 = n2876;
  assign po828 = n2877;
  assign po829 = n2878;
  assign po830 = n2879;
  assign po831 = n2880;
  assign po832 = n2881;
  assign po833 = n2882;
  assign po834 = n2883;
  assign po835 = n2884;
  assign po836 = n2885;
  assign po837 = n2886;
  assign po838 = n2887;
  assign po839 = n2888;
  assign po840 = n2889;
  assign po841 = n2890;
  assign po842 = n2891;
  assign po843 = n2892;
  assign po844 = n2893;
  assign po845 = n2894;
  assign po846 = n2895;
  assign po847 = n2896;
  assign po848 = n2897;
  assign po849 = n2898;
  assign po850 = n2899;
  assign po851 = n2900;
  assign po852 = n2901;
  assign po853 = n2902;
  assign po854 = n2903;
  assign po855 = n2904;
  assign po856 = n2905;
  assign po857 = n2906;
  assign po858 = n2907;
  assign po859 = n2908;
  assign po860 = n2909;
  assign po861 = n2910;
  assign po862 = n2911;
  assign po863 = n2912;
  assign po864 = n2913;
  assign po865 = n2914;
  assign po866 = n2915;
  assign po867 = n2916;
  assign po868 = n2917;
  assign po869 = n2918;
  assign po870 = n2919;
  assign po871 = n2920;
  assign po872 = n2921;
  assign po873 = n2922;
  assign po874 = n2923;
  assign po875 = n2924;
  assign po876 = n2925;
  assign po877 = n2926;
  assign po878 = n2927;
  assign po879 = n2928;
  assign po880 = n2929;
  assign po881 = n2930;
  assign po882 = n2931;
  assign po883 = n2932;
  assign po884 = n2933;
  assign po885 = n2934;
  assign po886 = n2935;
  assign po887 = n2936;
  assign po888 = n2937;
  assign po889 = n2938;
  assign po890 = n2939;
  assign po891 = n2940;
  assign po892 = n2941;
  assign po893 = n2942;
  assign po894 = n2943;
  assign po895 = n2944;
  assign po896 = n2945;
  assign po897 = n2946;
  assign po898 = n2947;
  assign po899 = n2948;
  assign po900 = n2949;
  assign po901 = n2950;
  assign po902 = n2951;
  assign po903 = n2952;
  assign po904 = n2953;
  assign po905 = n2954;
  assign po906 = n2955;
  assign po907 = n2956;
  assign po908 = n2957;
  assign po909 = n2958;
  assign po910 = n2959;
  assign po911 = n2960;
  assign po912 = n2961;
  assign po913 = n2962;
  assign po914 = n2963;
  assign po915 = n2964;
  assign po916 = n2965;
  assign po917 = n2966;
  assign po918 = n2967;
  assign po919 = n2968;
  assign po920 = n2969;
  assign po921 = n2970;
  assign po922 = n2971;
  assign po923 = n2972;
  assign po924 = n2973;
  assign po925 = n2974;
  assign po926 = n2975;
  assign po927 = n2976;
  assign po928 = n2977;
  assign po929 = n2978;
  assign po930 = n2979;
  assign po931 = n2980;
  assign po932 = n2981;
  assign po933 = n2982;
  assign po934 = n2983;
  assign po935 = n2984;
  assign po936 = n2985;
  assign po937 = n2986;
  assign po938 = n2987;
  assign po939 = n2988;
  assign po940 = n2989;
  assign po941 = n2990;
  assign po942 = n2991;
  assign po943 = n2992;
  assign po944 = n2993;
  assign po945 = n2994;
  assign po946 = n2995;
  assign po947 = n2996;
  assign po948 = n2997;
  assign po949 = n2998;
  assign po950 = n2999;
  assign po951 = n3000;
  assign po952 = n3001;
  assign po953 = n3002;
  assign po954 = n3003;
  assign po955 = n3004;
  assign po956 = n3005;
  assign po957 = n3006;
  assign po958 = n3007;
  assign po959 = n3008;
  assign po960 = n3009;
  assign po961 = n3010;
  assign po962 = n3011;
  assign po963 = n3012;
  assign po964 = n3013;
  assign po965 = n3014;
  assign po966 = n3015;
  assign po967 = n3016;
  assign po968 = n3017;
  assign po969 = n3018;
  assign po970 = n3019;
  assign po971 = n3020;
  assign po972 = n3021;
  assign po973 = n3022;
  assign po974 = n3023;
  assign po975 = n3024;
  assign po976 = n3025;
  assign po977 = n3026;
  assign po978 = n3027;
  assign po979 = n3028;
  assign po980 = n3029;
  assign po981 = n3030;
  assign po982 = n3031;
  assign po983 = n3032;
  assign po984 = n3033;
  assign po985 = n3034;
  assign po986 = n3035;
  assign po987 = n3036;
  assign po988 = n3037;
  assign po989 = n3038;
  assign po990 = n3039;
  assign po991 = n3040;
  assign po992 = n3041;
  assign po993 = n3042;
  assign po994 = n3043;
  assign po995 = n3044;
  assign po996 = n3045;
  assign po997 = n3046;
  assign po998 = n3047;
  assign po999 = n3048;
  assign po1000 = n3049;
  assign po1001 = n3050;
  assign po1002 = n3051;
  assign po1003 = n3052;
  assign po1004 = n3053;
  assign po1005 = n3054;
  assign po1006 = n3055;
  assign po1007 = n3056;
  assign po1008 = n3057;
  assign po1009 = n3058;
  assign po1010 = n3059;
  assign po1011 = n3060;
  assign po1012 = n3061;
  assign po1013 = n3062;
  assign po1014 = n3063;
  assign po1015 = n3064;
  assign po1016 = n3065;
  assign po1017 = n3066;
  assign po1018 = n3067;
  assign po1019 = n3068;
  assign po1020 = n3069;
  assign po1021 = n3070;
  assign po1022 = n3071;
  assign po1023 = n3072;
  assign po1024 = n3073;
  assign po1025 = n3074;
  assign po1026 = n3075;
  assign po1027 = n3076;
  assign po1028 = n3077;
  assign po1029 = n3078;
  assign po1030 = n3079;
  assign po1031 = n3080;
  assign po1032 = n3081;
  assign po1033 = n3082;
  assign po1034 = n3083;
  assign po1035 = n3084;
  assign po1036 = n3085;
  assign po1037 = n3086;
  assign po1038 = n3087;
  assign po1039 = n3088;
  assign po1040 = n3089;
  assign po1041 = n3090;
  assign po1042 = n3091;
  assign po1043 = n3092;
  assign po1044 = n3093;
  assign po1045 = n3094;
  assign po1046 = n3095;
  assign po1047 = n3096;
  assign po1048 = n3097;
  assign po1049 = n3098;
  assign po1050 = n3099;
  assign po1051 = n3100;
  assign po1052 = n3101;
  assign po1053 = n3102;
  assign po1054 = n3103;
  assign po1055 = n3104;
  assign po1056 = n3105;
  assign po1057 = n3106;
  assign po1058 = n3107;
  assign po1059 = n3108;
  assign po1060 = n3109;
  assign po1061 = n3110;
  assign po1062 = n3111;
  assign po1063 = n3112;
  assign po1064 = n3113;
  assign po1065 = n3114;
  assign po1066 = n3115;
  assign po1067 = n3116;
  assign po1068 = n3117;
  assign po1069 = n3118;
  assign po1070 = n3119;
  assign po1071 = n3120;
  assign po1072 = n3121;
  assign po1073 = n3122;
  assign po1074 = n3123;
  assign po1075 = n3124;
  assign po1076 = n3125;
  assign po1077 = n3126;
  assign po1078 = n3127;
  assign po1079 = n3128;
  assign po1080 = n3129;
  assign po1081 = n3130;
  assign po1082 = n3131;
  assign po1083 = n3132;
  assign po1084 = n3133;
  assign po1085 = n3134;
  assign po1086 = n3135;
  assign po1087 = n3136;
  assign po1088 = n3137;
  assign po1089 = n3138;
  assign po1090 = n3139;
  assign po1091 = n3140;
  assign po1092 = n3141;
  assign po1093 = n3142;
  assign po1094 = n3143;
  assign po1095 = n3144;
  assign po1096 = n3145;
  assign po1097 = n3146;
  assign po1098 = n3147;
  assign po1099 = n3148;
  assign po1100 = n3149;
  assign po1101 = n3150;
  assign po1102 = n3151;
  assign po1103 = n3152;
  assign po1104 = n3153;
  assign po1105 = n3154;
  assign po1106 = n3155;
  assign po1107 = n3156;
  assign po1108 = n3157;
  assign po1109 = n3158;
  assign po1110 = n3159;
  assign po1111 = n3160;
  assign po1112 = n3161;
  assign po1113 = n3162;
  assign po1114 = n3163;
  assign po1115 = n3164;
  assign po1116 = n3165;
  assign po1117 = n3166;
  assign po1118 = n3167;
  assign po1119 = n3168;
  assign po1120 = n3169;
  assign po1121 = n3170;
  assign po1122 = n3171;
  assign po1123 = n3172;
  assign po1124 = n3173;
  assign po1125 = n3174;
  assign po1126 = n3175;
  assign po1127 = n3176;
  assign po1128 = n3177;
  assign po1129 = n3178;
  assign po1130 = n3179;
  assign po1131 = n3180;
  assign po1132 = n3181;
  assign po1133 = n3182;
  assign po1134 = n3183;
  assign po1135 = n3184;
  assign po1136 = n3185;
  assign po1137 = n3186;
  assign po1138 = n3187;
  assign po1139 = n3188;
  assign po1140 = n3189;
  assign po1141 = n3190;
  assign po1142 = n3191;
  assign po1143 = n3192;
  assign po1144 = n3193;
  assign po1145 = n3194;
  assign po1146 = n3195;
  assign po1147 = n3196;
  assign po1148 = n3197;
  assign po1149 = n3198;
  assign po1150 = n3199;
  assign po1151 = n3200;
  assign po1152 = n3201;
  assign po1153 = n3202;
  assign po1154 = n3203;
  assign po1155 = n3204;
  assign po1156 = n3205;
  assign po1157 = n3206;
  assign po1158 = n3207;
  assign po1159 = n3208;
  assign po1160 = n3209;
  assign po1161 = n3210;
  assign po1162 = n3211;
  assign po1163 = n3212;
  assign po1164 = n3213;
  assign po1165 = n3214;
  assign po1166 = n3215;
  assign po1167 = n3216;
  assign po1168 = n3217;
  assign po1169 = n3218;
  assign po1170 = n3219;
  assign po1171 = n3220;
  assign po1172 = n3221;
  assign po1173 = n3222;
  assign po1174 = n3223;
  assign po1175 = n3224;
  assign po1176 = n3225;
  assign po1177 = n3226;
  assign po1178 = n3227;
  assign po1179 = n3228;
  assign po1180 = n3229;
  assign po1181 = n3230;
  assign po1182 = n3231;
  assign po1183 = n3232;
  assign po1184 = n3233;
  assign po1185 = n3234;
  assign po1186 = n3235;
  assign po1187 = n3236;
  assign po1188 = n3237;
  assign po1189 = n3238;
  assign po1190 = n3239;
  assign po1191 = n3240;
  assign po1192 = n3241;
  assign po1193 = n3242;
  assign po1194 = n3243;
  assign po1195 = n3244;
  assign po1196 = n3245;
  assign po1197 = n3246;
  assign po1198 = n3247;
  assign po1199 = n3248;
  assign po1200 = n3249;
  assign po1201 = n3250;
  assign po1202 = n3251;
  assign po1203 = n3252;
  assign po1204 = n3253;
  assign po1205 = n3254;
  assign po1206 = n3255;
  assign po1207 = n3256;
  assign po1208 = n3257;
  assign po1209 = n3258;
  assign po1210 = n3259;
  assign po1211 = n3260;
  assign po1212 = n3261;
  assign po1213 = n3262;
  assign po1214 = n3263;
  assign po1215 = n3264;
  assign po1216 = n3265;
  assign po1217 = n3266;
  assign po1218 = n3267;
  assign po1219 = n3268;
  assign po1220 = n3269;
  assign po1221 = n3270;
  assign po1222 = n3271;
  assign po1223 = n3272;
  assign po1224 = n3273;
  assign po1225 = n3274;
  assign po1226 = n3275;
  assign po1227 = n3276;
  assign po1228 = n3277;
  assign po1229 = n3278;
  assign po1230 = n3279;
  assign po1231 = n3280;
  assign po1232 = n3281;
  assign po1233 = n3282;
  assign po1234 = n3283;
  assign po1235 = n3284;
  assign po1236 = n3285;
  assign po1237 = n3286;
  assign po1238 = n3287;
  assign po1239 = n3288;
  assign po1240 = n3289;
  assign po1241 = n3290;
  assign po1242 = n3291;
  assign po1243 = n3292;
  assign po1244 = n3293;
  assign po1245 = n3294;
  assign po1246 = n3295;
  assign po1247 = n3296;
  assign po1248 = n3297;
  assign po1249 = n3298;
  assign po1250 = n3299;
  assign po1251 = n3300;
  assign po1252 = n3301;
  assign po1253 = n3302;
  assign po1254 = n3303;
  assign po1255 = n3304;
  assign po1256 = n3305;
  assign po1257 = n3306;
  assign po1258 = n3307;
  assign po1259 = n3308;
  assign po1260 = n3309;
  assign po1261 = n3310;
  assign po1262 = n3311;
  assign po1263 = n3312;
  assign po1264 = n3313;
  assign po1265 = n3314;
  assign po1266 = n3315;
  assign po1267 = n3316;
  assign po1268 = n3317;
  assign po1269 = n3318;
  assign po1270 = n3319;
  assign po1271 = n3320;
  assign po1272 = n3321;
  assign po1273 = n3322;
  assign po1274 = n3323;
  assign po1275 = n3324;
  assign po1276 = n3325;
  assign po1277 = n3326;
  assign po1278 = n3327;
  assign po1279 = n3328;
  assign po1280 = n3329;
  assign po1281 = n3330;
  assign po1282 = n3331;
  assign po1283 = n3332;
  assign po1284 = n3333;
  assign po1285 = n3334;
  assign po1286 = n3335;
  assign po1287 = n3336;
  assign po1288 = n3337;
  assign po1289 = n3338;
  assign po1290 = n3339;
  assign po1291 = n3340;
  assign po1292 = n3341;
  assign po1293 = n3342;
  assign po1294 = n3343;
  assign po1295 = n3344;
  assign po1296 = n3345;
  assign po1297 = n3346;
  assign po1298 = n3347;
  assign po1299 = n3348;
  assign po1300 = n3349;
  assign po1301 = n3350;
  assign po1302 = n3351;
  assign po1303 = n3352;
  assign po1304 = n3353;
  assign po1305 = n3354;
  assign po1306 = n3355;
  assign po1307 = n3356;
  assign po1308 = n3357;
  assign po1309 = n3358;
  assign po1310 = n3359;
  assign po1311 = n3360;
  assign po1312 = n3361;
  assign po1313 = n3362;
  assign po1314 = n3363;
  assign po1315 = n3364;
  assign po1316 = n3365;
  assign po1317 = n3366;
  assign po1318 = n3367;
  assign po1319 = n3368;
  assign po1320 = n3369;
  assign po1321 = n3370;
  assign po1322 = n3371;
  assign po1323 = n3372;
  assign po1324 = n3373;
  assign po1325 = n3374;
  assign po1326 = n3375;
  assign po1327 = n3376;
  assign po1328 = n3377;
  assign po1329 = n3378;
  assign po1330 = n3379;
  assign po1331 = n3380;
  assign po1332 = n3381;
  assign po1333 = n3382;
  assign po1334 = n3383;
  assign po1335 = n3384;
  assign po1336 = n3385;
  assign po1337 = n3386;
  assign po1338 = n3387;
  assign po1339 = n3388;
  assign po1340 = n3389;
  assign po1341 = n3390;
  assign po1342 = n3391;
  assign po1343 = n3392;
  assign po1344 = n3393;
  assign po1345 = n3394;
  assign po1346 = n3395;
  assign po1347 = n3396;
  assign po1348 = n3397;
  assign po1349 = n3398;
  assign po1350 = n3399;
  assign po1351 = n3400;
  assign po1352 = n3401;
  assign po1353 = n3402;
  assign po1354 = n3403;
  assign po1355 = n3404;
  assign po1356 = n3405;
  assign po1357 = n3406;
  assign po1358 = n3407;
  assign po1359 = n3408;
  assign po1360 = n3409;
  assign po1361 = n3410;
  assign po1362 = n3411;
  assign po1363 = n3412;
  assign po1364 = n3413;
  assign po1365 = n3414;
  assign po1366 = n3415;
  assign po1367 = n3416;
  assign po1368 = n3417;
  assign po1369 = n3418;
  assign po1370 = n3419;
  assign po1371 = n3420;
  assign po1372 = n3421;
  assign po1373 = n3422;
  assign po1374 = n3423;
  assign po1375 = n3424;
  assign po1376 = n3425;
  assign po1377 = n3426;
  assign po1378 = n3427;
  assign po1379 = n3428;
  assign po1380 = n3429;
  assign po1381 = n3430;
  assign po1382 = n3431;
  assign po1383 = n3432;
  assign po1384 = n3433;
  assign po1385 = n3434;
  assign po1386 = n3435;
  assign po1387 = n3436;
  assign po1388 = n3437;
  assign po1389 = n3438;
  assign po1390 = n3439;
  assign po1391 = n3440;
  assign po1392 = n3441;
  assign po1393 = n3442;
  assign po1394 = n3443;
  assign po1395 = n3444;
  assign po1396 = n3445;
  assign po1397 = n3446;
  assign po1398 = n3447;
  assign po1399 = n3448;
  assign po1400 = n3449;
  assign po1401 = n3450;
  assign po1402 = n3451;
  assign po1403 = n3452;
  assign po1404 = n3453;
  assign po1405 = n3454;
  assign po1406 = n3455;
  assign po1407 = n3456;
  assign po1408 = n3457;
  assign po1409 = n3458;
  assign po1410 = n3459;
  assign po1411 = n3460;
  assign po1412 = n3461;
  assign po1413 = n3462;
  assign po1414 = n3463;
  assign po1415 = n3464;
  assign po1416 = n3465;
  assign po1417 = n3466;
  assign po1418 = n3467;
  assign po1419 = n3468;
  assign po1420 = n3469;
  assign po1421 = n3470;
  assign po1422 = n3471;
  assign po1423 = n3472;
  assign po1424 = n3473;
  assign po1425 = n3474;
  assign po1426 = n3475;
  assign po1427 = n3476;
  assign po1428 = n3477;
  assign po1429 = n3478;
  assign po1430 = n3479;
  assign po1431 = n3480;
  assign po1432 = n3481;
  assign po1433 = n3482;
  assign po1434 = n3483;
  assign po1435 = n3484;
  assign po1436 = n3485;
  assign po1437 = n3486;
  assign po1438 = n3487;
  assign po1439 = n3488;
  assign po1440 = n3489;
  assign po1441 = n3490;
  assign po1442 = n3491;
  assign po1443 = n3492;
  assign po1444 = n3493;
  assign po1445 = n3494;
  assign po1446 = n3495;
  assign po1447 = n3496;
  assign po1448 = n3497;
  assign po1449 = n3498;
  assign po1450 = n3499;
  assign po1451 = n3500;
  assign po1452 = n3501;
  assign po1453 = n3502;
  assign po1454 = n3503;
  assign po1455 = n3504;
  assign po1456 = n3505;
  assign po1457 = n3506;
  assign po1458 = n3507;
  assign po1459 = n3508;
  assign po1460 = n3509;
  assign po1461 = n3510;
  assign po1462 = n3511;
  assign po1463 = n3512;
  assign po1464 = n3513;
  assign po1465 = n3514;
  assign po1466 = n3515;
  assign po1467 = n3516;
  assign po1468 = n3517;
  assign po1469 = n3518;
  assign po1470 = n3519;
  assign po1471 = n3520;
  assign po1472 = n3521;
  assign po1473 = n3522;
  assign po1474 = n3523;
  assign po1475 = n3524;
  assign po1476 = n3525;
  assign po1477 = n3526;
  assign po1478 = n3527;
  assign po1479 = n3528;
  assign po1480 = n3529;
  assign po1481 = n3530;
  assign po1482 = n3531;
  assign po1483 = n3532;
  assign po1484 = n3533;
  assign po1485 = n3534;
  assign po1486 = n3535;
  assign po1487 = n3536;
  assign po1488 = n3537;
  assign po1489 = n3538;
  assign po1490 = n3539;
  assign po1491 = n3540;
  assign po1492 = n3541;
  assign po1493 = n3542;
  assign po1494 = n3543;
  assign po1495 = n3544;
  assign po1496 = n3545;
  assign po1497 = n3546;
  assign po1498 = n3547;
  assign po1499 = n3548;
  assign po1500 = n3549;
  assign po1501 = n3550;
  assign po1502 = n3551;
  assign po1503 = n3552;
  assign po1504 = n3553;
  assign po1505 = n3554;
  assign po1506 = n3555;
  assign po1507 = n3556;
  assign po1508 = n3557;
  assign po1509 = n3558;
  assign po1510 = n3559;
  assign po1511 = n3560;
  assign po1512 = n3561;
  assign po1513 = n3562;
  assign po1514 = n3563;
  assign po1515 = n3564;
  assign po1516 = n3565;
  assign po1517 = n3566;
  assign po1518 = n3567;
  assign po1519 = n3568;
  assign po1520 = n3569;
  assign po1521 = n3570;
  assign po1522 = n3571;
  assign po1523 = n3572;
  assign po1524 = n3573;
  assign po1525 = n3574;
  assign po1526 = n3575;
  assign po1527 = n3576;
  assign po1528 = n3577;
  assign po1529 = n3578;
  assign po1530 = n3579;
  assign po1531 = n3580;
  assign po1532 = n3581;
  assign po1533 = n3582;
  assign po1534 = n3583;
  assign po1535 = n3584;
  assign po1536 = n3585;
  assign po1537 = n3586;
  assign po1538 = n3587;
  assign po1539 = n3588;
  assign po1540 = n3589;
  assign po1541 = n3590;
  assign po1542 = n3591;
  assign po1543 = n3592;
  assign po1544 = n3593;
  assign po1545 = n3594;
  assign po1546 = n3595;
  assign po1547 = n3596;
  assign po1548 = n3597;
  assign po1549 = n3598;
  assign po1550 = n3599;
  assign po1551 = n3600;
  assign po1552 = n3601;
  assign po1553 = n3602;
  assign po1554 = n3603;
  assign po1555 = n3604;
  assign po1556 = n3605;
  assign po1557 = n3606;
  assign po1558 = n3607;
  assign po1559 = n3608;
  assign po1560 = n3609;
  assign po1561 = n3610;
  assign po1562 = n3611;
  assign po1563 = n3612;
  assign po1564 = n3613;
  assign po1565 = n3614;
  assign po1566 = n3615;
  assign po1567 = n3616;
  assign po1568 = n3617;
  assign po1569 = n3618;
  assign po1570 = n3619;
  assign po1571 = n3620;
  assign po1572 = n3621;
  assign po1573 = n3622;
  assign po1574 = n3623;
  assign po1575 = n3624;
  assign po1576 = n3625;
  assign po1577 = n3626;
  assign po1578 = n3627;
  assign po1579 = n3628;
  assign po1580 = n3629;
  assign po1581 = n3630;
  assign po1582 = n3631;
  assign po1583 = n3632;
  assign po1584 = n3633;
  assign po1585 = n3634;
  assign po1586 = n3635;
  assign po1587 = n3636;
  assign po1588 = n3637;
  assign po1589 = n3638;
  assign po1590 = n3639;
  assign po1591 = n3640;
  assign po1592 = n3641;
  assign po1593 = n3642;
  assign po1594 = n3643;
  assign po1595 = n3644;
  assign po1596 = n3645;
  assign po1597 = n3646;
  assign po1598 = n3647;
  assign po1599 = n3648;
  assign po1600 = n3649;
  assign po1601 = n3650;
  assign po1602 = n3651;
  assign po1603 = n3652;
  assign po1604 = n3653;
  assign po1605 = n3654;
  assign po1606 = n3655;
  assign po1607 = n3656;
  assign po1608 = n3657;
  assign po1609 = n3658;
  assign po1610 = n3659;
  assign po1611 = n3660;
  assign po1612 = n3661;
  assign po1613 = n3662;
  assign po1614 = n3663;
  assign po1615 = n3664;
  assign po1616 = n3665;
  assign po1617 = n3666;
  assign po1618 = n3667;
  assign po1619 = n3668;
  assign po1620 = n3669;
  assign po1621 = n3670;
  assign po1622 = n3671;
  assign po1623 = n3672;
  assign po1624 = n3673;
  assign po1625 = n3674;
  assign po1626 = n3675;
  assign po1627 = n3676;
  assign po1628 = n3677;
  assign po1629 = n3678;
  assign po1630 = n3679;
  assign po1631 = n3680;
  assign po1632 = n3681;
  assign po1633 = n3682;
  assign po1634 = n3683;
  assign po1635 = n3684;
  assign po1636 = n3685;
  assign po1637 = n3686;
  assign po1638 = n3687;
  assign po1639 = n3688;
  assign po1640 = n3689;
  assign po1641 = n3690;
  assign po1642 = n3691;
  assign po1643 = n3692;
  assign po1644 = n3693;
  assign po1645 = n3694;
  assign po1646 = n3695;
  assign po1647 = n3696;
  assign po1648 = n3697;
  assign po1649 = n3698;
  assign po1650 = n3699;
  assign po1651 = n3700;
  assign po1652 = n3701;
  assign po1653 = n3702;
  assign po1654 = n3703;
  assign po1655 = n3704;
  assign po1656 = n3705;
  assign po1657 = n3706;
  assign po1658 = n3707;
  assign po1659 = n3708;
  assign po1660 = n3709;
  assign po1661 = n3710;
  assign po1662 = n3711;
  assign po1663 = n3712;
  assign po1664 = n3713;
  assign po1665 = n3714;
  assign po1666 = n3715;
  assign po1667 = n3716;
  assign po1668 = n3717;
  assign po1669 = n3718;
  assign po1670 = n3719;
  assign po1671 = n3720;
  assign po1672 = n3721;
  assign po1673 = n3722;
  assign po1674 = n3723;
  assign po1675 = n3724;
  assign po1676 = n3725;
  assign po1677 = n3726;
  assign po1678 = n3727;
  assign po1679 = n3728;
  assign po1680 = n3729;
  assign po1681 = n3730;
  assign po1682 = n3731;
  assign po1683 = n3732;
  assign po1684 = n3733;
  assign po1685 = n3734;
  assign po1686 = n3735;
  assign po1687 = n3736;
  assign po1688 = n3737;
  assign po1689 = n3738;
  assign po1690 = n3739;
  assign po1691 = n3740;
  assign po1692 = n3741;
  assign po1693 = n3742;
  assign po1694 = n3743;
  assign po1695 = n3744;
  assign po1696 = n3745;
  assign po1697 = n3746;
  assign po1698 = n3747;
  assign po1699 = n3748;
  assign po1700 = n3749;
  assign po1701 = n3750;
  assign po1702 = n3751;
  assign po1703 = n3752;
  assign po1704 = n3753;
  assign po1705 = n3754;
  assign po1706 = n3755;
  assign po1707 = n3756;
  assign po1708 = n3757;
  assign po1709 = n3758;
  assign po1710 = n3759;
  assign po1711 = n3760;
  assign po1712 = n3761;
  assign po1713 = n3762;
  assign po1714 = n3763;
  assign po1715 = n3764;
  assign po1716 = n3765;
  assign po1717 = n3766;
  assign po1718 = n3767;
  assign po1719 = n3768;
  assign po1720 = n3769;
  assign po1721 = n3770;
  assign po1722 = n3771;
  assign po1723 = n3772;
  assign po1724 = n3773;
  assign po1725 = n3774;
  assign po1726 = n3775;
  assign po1727 = n3776;
  assign po1728 = n3777;
  assign po1729 = n3778;
  assign po1730 = n3779;
  assign po1731 = n3780;
  assign po1732 = n3781;
  assign po1733 = n3782;
  assign po1734 = n3783;
  assign po1735 = n3784;
  assign po1736 = n3785;
  assign po1737 = n3786;
  assign po1738 = n3787;
  assign po1739 = n3788;
  assign po1740 = n3789;
  assign po1741 = n3790;
  assign po1742 = n3791;
  assign po1743 = n3792;
  assign po1744 = n3793;
  assign po1745 = n3794;
  assign po1746 = n3795;
  assign po1747 = n3796;
  assign po1748 = n3797;
  assign po1749 = n3798;
  assign po1750 = n3799;
  assign po1751 = n3800;
  assign po1752 = n3801;
  assign po1753 = n3802;
  assign po1754 = n3803;
  assign po1755 = n3804;
  assign po1756 = n3805;
  assign po1757 = n3806;
  assign po1758 = n3807;
  assign po1759 = n3808;
  assign po1760 = n3809;
  assign po1761 = n3810;
  assign po1762 = n3811;
  assign po1763 = n3812;
  assign po1764 = n3813;
  assign po1765 = n3814;
  assign po1766 = n3815;
  assign po1767 = n3816;
  assign po1768 = n3817;
  assign po1769 = n3818;
  assign po1770 = n3819;
  assign po1771 = n3820;
  assign po1772 = n3821;
  assign po1773 = n3822;
  assign po1774 = n3823;
  assign po1775 = n3824;
  assign po1776 = n3825;
  assign po1777 = n3826;
  assign po1778 = n3827;
  assign po1779 = n3828;
  assign po1780 = n3829;
  assign po1781 = n3830;
  assign po1782 = n3831;
  assign po1783 = n3832;
  assign po1784 = n3833;
  assign po1785 = n3834;
  assign po1786 = n3835;
  assign po1787 = n3836;
  assign po1788 = n3837;
  assign po1789 = n3838;
  assign po1790 = n3839;
  assign po1791 = n3840;
  assign po1792 = n3841;
  assign po1793 = n3842;
  assign po1794 = n3843;
  assign po1795 = n3844;
  assign po1796 = n3845;
  assign po1797 = n3846;
  assign po1798 = n3847;
  assign po1799 = n3848;
  assign po1800 = n3849;
  assign po1801 = n3850;
  assign po1802 = n3851;
  assign po1803 = n3852;
  assign po1804 = n3853;
  assign po1805 = n3854;
  assign po1806 = n3855;
  assign po1807 = n3856;
  assign po1808 = n3857;
  assign po1809 = n3858;
  assign po1810 = n3859;
  assign po1811 = n3860;
  assign po1812 = n3861;
  assign po1813 = n3862;
  assign po1814 = n3863;
  assign po1815 = n3864;
  assign po1816 = n3865;
  assign po1817 = n3866;
  assign po1818 = n3867;
  assign po1819 = n3868;
  assign po1820 = n3869;
  assign po1821 = n3870;
  assign po1822 = n3871;
  assign po1823 = n3872;
  assign po1824 = n3873;
  assign po1825 = n3874;
  assign po1826 = n3875;
  assign po1827 = n3876;
  assign po1828 = n3877;
  assign po1829 = n3878;
  assign po1830 = n3879;
  assign po1831 = n3880;
  assign po1832 = n3881;
  assign po1833 = n3882;
  assign po1834 = n3883;
  assign po1835 = n3884;
  assign po1836 = n3885;
  assign po1837 = n3886;
  assign po1838 = n3887;
  assign po1839 = n3888;
  assign po1840 = n3889;
  assign po1841 = n3890;
  assign po1842 = n3891;
  assign po1843 = n3892;
  assign po1844 = n3893;
  assign po1845 = n3894;
  assign po1846 = n3895;
  assign po1847 = n3896;
  assign po1848 = n3897;
  assign po1849 = n3898;
  assign po1850 = n3899;
  assign po1851 = n3900;
  assign po1852 = n3901;
  assign po1853 = n3902;
  assign po1854 = n3903;
  assign po1855 = n3904;
  assign po1856 = n3905;
  assign po1857 = n3906;
  assign po1858 = n3907;
  assign po1859 = n3908;
  assign po1860 = n3909;
  assign po1861 = n3910;
  assign po1862 = n3911;
  assign po1863 = n3912;
  assign po1864 = n3913;
  assign po1865 = n3914;
  assign po1866 = n3915;
  assign po1867 = n3916;
  assign po1868 = n3917;
  assign po1869 = n3918;
  assign po1870 = n3919;
  assign po1871 = n3920;
  assign po1872 = n3921;
  assign po1873 = n3922;
  assign po1874 = n3923;
  assign po1875 = n3924;
  assign po1876 = n3925;
  assign po1877 = n3926;
  assign po1878 = n3927;
  assign po1879 = n3928;
  assign po1880 = n3929;
  assign po1881 = n3930;
  assign po1882 = n3931;
  assign po1883 = n3932;
  assign po1884 = n3933;
  assign po1885 = n3934;
  assign po1886 = n3935;
  assign po1887 = n3936;
  assign po1888 = n3937;
  assign po1889 = n3938;
  assign po1890 = n3939;
  assign po1891 = n3940;
  assign po1892 = n3941;
  assign po1893 = n3942;
  assign po1894 = n3943;
  assign po1895 = n3944;
  assign po1896 = n3945;
  assign po1897 = n3946;
  assign po1898 = n3947;
  assign po1899 = n3948;
  assign po1900 = n3949;
  assign po1901 = n3950;
  assign po1902 = n3951;
  assign po1903 = n3952;
  assign po1904 = n3953;
  assign po1905 = n3954;
  assign po1906 = n3955;
  assign po1907 = n3956;
  assign po1908 = n3957;
  assign po1909 = n3958;
  assign po1910 = n3959;
  assign po1911 = n3960;
  assign po1912 = n3961;
  assign po1913 = n3962;
  assign po1914 = n3963;
  assign po1915 = n3964;
  assign po1916 = n3965;
  assign po1917 = n3966;
  assign po1918 = n3967;
  assign po1919 = n3968;
  assign po1920 = n3969;
  assign po1921 = n3970;
  assign po1922 = n3971;
  assign po1923 = n3972;
  assign po1924 = n3973;
  assign po1925 = n3974;
  assign po1926 = n3975;
  assign po1927 = n3976;
  assign po1928 = n3977;
  assign po1929 = n3978;
  assign po1930 = n3979;
  assign po1931 = n3980;
  assign po1932 = n3981;
  assign po1933 = n3982;
  assign po1934 = n3983;
  assign po1935 = n3984;
  assign po1936 = n3985;
  assign po1937 = n3986;
  assign po1938 = n3987;
  assign po1939 = n3988;
  assign po1940 = n3989;
  assign po1941 = n3990;
  assign po1942 = n3991;
  assign po1943 = n3992;
  assign po1944 = n3993;
  assign po1945 = n3994;
  assign po1946 = n3995;
  assign po1947 = n3996;
  assign po1948 = n3997;
  assign po1949 = n3998;
  assign po1950 = n3999;
  assign po1951 = n4000;
  assign po1952 = n4001;
  assign po1953 = n4002;
  assign po1954 = n4003;
  assign po1955 = n4004;
  assign po1956 = n4005;
  assign po1957 = n4006;
  assign po1958 = n4007;
  assign po1959 = n4008;
  assign po1960 = n4009;
  assign po1961 = n4010;
  assign po1962 = n4011;
  assign po1963 = n4012;
  assign po1964 = n4013;
  assign po1965 = n4014;
  assign po1966 = n4015;
  assign po1967 = n4016;
  assign po1968 = n4017;
  assign po1969 = n4018;
  assign po1970 = n4019;
  assign po1971 = n4020;
  assign po1972 = n4021;
  assign po1973 = n4022;
  assign po1974 = n4023;
  assign po1975 = n4024;
  assign po1976 = n4025;
  assign po1977 = n4026;
  assign po1978 = n4027;
  assign po1979 = n4028;
  assign po1980 = n4029;
  assign po1981 = n4030;
  assign po1982 = n4031;
  assign po1983 = n4032;
  assign po1984 = n4033;
  assign po1985 = n4034;
  assign po1986 = n4035;
  assign po1987 = n4036;
  assign po1988 = n4037;
  assign po1989 = n4038;
  assign po1990 = n4039;
  assign po1991 = n4040;
  assign po1992 = n4041;
  assign po1993 = n4042;
  assign po1994 = n4043;
  assign po1995 = n4044;
  assign po1996 = n4045;
  assign po1997 = n4046;
  assign po1998 = n4047;
  assign po1999 = n4048;
  assign po2000 = n4049;
  assign po2001 = n4050;
  assign po2002 = n4051;
  assign po2003 = n4052;
  assign po2004 = n4053;
  assign po2005 = n4054;
  assign po2006 = n4055;
  assign po2007 = n4056;
  assign po2008 = n4057;
  assign po2009 = n4058;
  assign po2010 = n4059;
  assign po2011 = n4060;
  assign po2012 = n4061;
  assign po2013 = n4062;
  assign po2014 = n4063;
  assign po2015 = n4064;
  assign po2016 = n4065;
  assign po2017 = n4066;
  assign po2018 = n4067;
  assign po2019 = n4068;
  assign po2020 = n4069;
  assign po2021 = n4070;
  assign po2022 = n4071;
  assign po2023 = n4072;
  assign po2024 = n4073;
  assign po2025 = n4074;
  assign po2026 = n4075;
  assign po2027 = n4076;
  assign po2028 = n4077;
  assign po2029 = n4078;
  assign po2030 = n4079;
  assign po2031 = n4080;
  assign po2032 = n4081;
  assign po2033 = n4082;
  assign po2034 = n4083;
  assign po2035 = n4084;
  assign po2036 = n4085;
  assign po2037 = n4086;
  assign po2038 = n4087;
  assign po2039 = n4088;
  assign po2040 = n4089;
  assign po2041 = n4090;
  assign po2042 = n4091;
  assign po2043 = n4092;
  assign po2044 = n4093;
  assign po2045 = n4094;
  assign po2046 = n4095;
  assign po2047 = n4096;
  assign po2048 = ~new_n5280;
  assign po2049 = ~new_n5282;
  assign po2050 = ~new_n5284;
  assign po2051 = ~new_n5288;
  assign po2052 = ~new_n5292;
  assign po2053 = ~new_n5296;
  assign po2054 = ~new_n5300;
  assign po2055 = ~new_n5304;
  assign po2056 = ~new_n5308;
  assign po2057 = ~new_n5312;
  assign po2058 = ~new_n5316;
  assign po2059 = ~new_n5320;
  assign po2060 = ~new_n5324;
  assign po2061 = ~new_n5328;
  assign po2062 = ~new_n5334;
  assign po2063 = ~new_n5340;
  assign po2064 = ~new_n5346;
  assign po2065 = ~new_n5352;
  assign po2066 = ~new_n5358;
  assign po2067 = ~new_n5364;
  assign po2068 = ~new_n5370;
  assign po2069 = ~new_n5376;
  assign po2070 = ~new_n5382;
  assign po2071 = ~new_n5388;
  assign po2072 = ~new_n5394;
  assign po2073 = ~new_n5400;
  assign po2074 = ~new_n5406;
  assign po2075 = ~new_n5412;
  assign po2076 = ~new_n5414;
  assign po2077 = ~new_n5421;
  assign po2078 = n32;
  assign po2079 = n31;
  assign po2080 = n30;
  assign po2081 = n29;
  assign po2082 = n28;
  assign po2083 = n27;
  assign po2084 = n26;
  assign po2085 = n25;
  assign po2086 = n24;
  assign po2087 = n23;
  assign po2088 = n22;
  assign po2089 = n21;
  assign po2090 = n20;
  assign po2091 = n19;
  assign po2092 = n18;
  assign po2093 = n17;
  assign po2094 = n16;
  assign po2095 = n15;
  assign po2096 = n14;
  assign po2097 = n13;
  assign po2098 = n12;
  assign po2099 = n11;
  assign po2100 = n10;
  assign po2101 = n9;
  assign po2102 = n8;
  assign po2103 = n7;
  assign po2104 = n6;
  assign po2105 = n5;
  assign po2106 = n4;
  assign po2107 = n3;
  assign po2108 = n2;
  assign po2109 = n1;
  assign po2110 = n64;
  assign po2111 = n63;
  assign po2112 = n62;
  assign po2113 = n61;
  assign po2114 = n60;
  assign po2115 = n59;
  assign po2116 = n58;
  assign po2117 = n57;
  assign po2118 = n56;
  assign po2119 = n55;
  assign po2120 = n54;
  assign po2121 = n53;
  assign po2122 = n52;
  assign po2123 = n51;
  assign po2124 = n50;
  assign po2125 = n49;
  assign po2126 = n48;
  assign po2127 = n47;
  assign po2128 = n46;
  assign po2129 = n45;
  assign po2130 = n44;
  assign po2131 = n43;
  assign po2132 = n42;
  assign po2133 = n41;
  assign po2134 = n40;
  assign po2135 = n39;
  assign po2136 = n38;
  assign po2137 = n37;
  assign po2138 = n36;
  assign po2139 = n35;
  assign po2140 = n34;
  assign po2141 = n33;
  assign po2142 = n96;
  assign po2143 = n95;
  assign po2144 = n94;
  assign po2145 = n93;
  assign po2146 = n92;
  assign po2147 = n91;
  assign po2148 = n90;
  assign po2149 = n89;
  assign po2150 = n88;
  assign po2151 = n87;
  assign po2152 = n86;
  assign po2153 = n85;
  assign po2154 = n84;
  assign po2155 = n83;
  assign po2156 = n82;
  assign po2157 = n81;
  assign po2158 = n80;
  assign po2159 = n79;
  assign po2160 = n78;
  assign po2161 = n77;
  assign po2162 = n76;
  assign po2163 = n75;
  assign po2164 = n74;
  assign po2165 = n73;
  assign po2166 = n72;
  assign po2167 = n71;
  assign po2168 = n70;
  assign po2169 = n69;
  assign po2170 = n68;
  assign po2171 = n67;
  assign po2172 = n66;
  assign po2173 = n65;
  assign po2174 = n128;
  assign po2175 = n127;
  assign po2176 = n126;
  assign po2177 = n125;
  assign po2178 = n124;
  assign po2179 = n123;
  assign po2180 = n122;
  assign po2181 = n121;
  assign po2182 = n120;
  assign po2183 = n119;
  assign po2184 = n118;
  assign po2185 = n117;
  assign po2186 = n116;
  assign po2187 = n115;
  assign po2188 = n114;
  assign po2189 = n113;
  assign po2190 = n112;
  assign po2191 = n111;
  assign po2192 = n110;
  assign po2193 = n109;
  assign po2194 = n108;
  assign po2195 = n107;
  assign po2196 = n106;
  assign po2197 = n105;
  assign po2198 = n104;
  assign po2199 = n103;
  assign po2200 = n102;
  assign po2201 = n101;
  assign po2202 = n100;
  assign po2203 = n99;
  assign po2204 = n98;
  assign po2205 = n97;
  assign po2206 = n160;
  assign po2207 = n159;
  assign po2208 = n158;
  assign po2209 = n157;
  assign po2210 = n156;
  assign po2211 = n155;
  assign po2212 = n154;
  assign po2213 = n153;
  assign po2214 = n152;
  assign po2215 = n151;
  assign po2216 = n150;
  assign po2217 = n149;
  assign po2218 = n148;
  assign po2219 = n147;
  assign po2220 = n146;
  assign po2221 = n145;
  assign po2222 = n144;
  assign po2223 = n143;
  assign po2224 = n142;
  assign po2225 = n141;
  assign po2226 = n140;
  assign po2227 = n139;
  assign po2228 = n138;
  assign po2229 = n137;
  assign po2230 = n136;
  assign po2231 = n135;
  assign po2232 = n134;
  assign po2233 = n133;
  assign po2234 = n132;
  assign po2235 = n131;
  assign po2236 = n130;
  assign po2237 = n129;
  assign po2238 = n192;
  assign po2239 = n191;
  assign po2240 = n190;
  assign po2241 = n189;
  assign po2242 = n188;
  assign po2243 = n187;
  assign po2244 = n186;
  assign po2245 = n185;
  assign po2246 = n184;
  assign po2247 = n183;
  assign po2248 = n182;
  assign po2249 = n181;
  assign po2250 = n180;
  assign po2251 = n179;
  assign po2252 = n178;
  assign po2253 = n177;
  assign po2254 = n176;
  assign po2255 = n175;
  assign po2256 = n174;
  assign po2257 = n173;
  assign po2258 = n172;
  assign po2259 = n171;
  assign po2260 = n170;
  assign po2261 = n169;
  assign po2262 = n168;
  assign po2263 = n167;
  assign po2264 = n166;
  assign po2265 = n165;
  assign po2266 = n164;
  assign po2267 = n163;
  assign po2268 = n162;
  assign po2269 = n161;
  assign po2270 = n224;
  assign po2271 = n223;
  assign po2272 = n222;
  assign po2273 = n221;
  assign po2274 = n220;
  assign po2275 = n219;
  assign po2276 = n218;
  assign po2277 = n217;
  assign po2278 = n216;
  assign po2279 = n215;
  assign po2280 = n214;
  assign po2281 = n213;
  assign po2282 = n212;
  assign po2283 = n211;
  assign po2284 = n210;
  assign po2285 = n209;
  assign po2286 = n208;
  assign po2287 = n207;
  assign po2288 = n206;
  assign po2289 = n205;
  assign po2290 = n204;
  assign po2291 = n203;
  assign po2292 = n202;
  assign po2293 = n201;
  assign po2294 = n200;
  assign po2295 = n199;
  assign po2296 = n198;
  assign po2297 = n197;
  assign po2298 = n196;
  assign po2299 = n195;
  assign po2300 = n194;
  assign po2301 = n193;
  assign po2302 = n256;
  assign po2303 = n255;
  assign po2304 = n254;
  assign po2305 = n253;
  assign po2306 = n252;
  assign po2307 = n251;
  assign po2308 = n250;
  assign po2309 = n249;
  assign po2310 = n248;
  assign po2311 = n247;
  assign po2312 = n246;
  assign po2313 = n245;
  assign po2314 = n244;
  assign po2315 = n243;
  assign po2316 = n242;
  assign po2317 = n241;
  assign po2318 = n240;
  assign po2319 = n239;
  assign po2320 = n238;
  assign po2321 = n237;
  assign po2322 = n236;
  assign po2323 = n235;
  assign po2324 = n234;
  assign po2325 = n233;
  assign po2326 = n232;
  assign po2327 = n231;
  assign po2328 = n230;
  assign po2329 = n229;
  assign po2330 = n228;
  assign po2331 = n227;
  assign po2332 = n226;
  assign po2333 = n225;
  assign po2334 = n288;
  assign po2335 = n287;
  assign po2336 = n286;
  assign po2337 = n285;
  assign po2338 = n284;
  assign po2339 = n283;
  assign po2340 = n282;
  assign po2341 = n281;
  assign po2342 = n280;
  assign po2343 = n279;
  assign po2344 = n278;
  assign po2345 = n277;
  assign po2346 = n276;
  assign po2347 = n275;
  assign po2348 = n274;
  assign po2349 = n273;
  assign po2350 = n272;
  assign po2351 = n271;
  assign po2352 = n270;
  assign po2353 = n269;
  assign po2354 = n268;
  assign po2355 = n267;
  assign po2356 = n266;
  assign po2357 = n265;
  assign po2358 = n264;
  assign po2359 = n263;
  assign po2360 = n262;
  assign po2361 = n261;
  assign po2362 = n260;
  assign po2363 = n259;
  assign po2364 = n258;
  assign po2365 = n257;
  assign po2366 = n320;
  assign po2367 = n319;
  assign po2368 = n318;
  assign po2369 = n317;
  assign po2370 = n316;
  assign po2371 = n315;
  assign po2372 = n314;
  assign po2373 = n313;
  assign po2374 = n312;
  assign po2375 = n311;
  assign po2376 = n310;
  assign po2377 = n309;
  assign po2378 = n308;
  assign po2379 = n307;
  assign po2380 = n306;
  assign po2381 = n305;
  assign po2382 = n304;
  assign po2383 = n303;
  assign po2384 = n302;
  assign po2385 = n301;
  assign po2386 = n300;
  assign po2387 = n299;
  assign po2388 = n298;
  assign po2389 = n297;
  assign po2390 = n296;
  assign po2391 = n295;
  assign po2392 = n294;
  assign po2393 = n293;
  assign po2394 = n292;
  assign po2395 = n291;
  assign po2396 = n290;
  assign po2397 = n289;
  assign po2398 = n352;
  assign po2399 = n351;
  assign po2400 = n350;
  assign po2401 = n349;
  assign po2402 = n348;
  assign po2403 = n347;
  assign po2404 = n346;
  assign po2405 = n345;
  assign po2406 = n344;
  assign po2407 = n343;
  assign po2408 = n342;
  assign po2409 = n341;
  assign po2410 = n340;
  assign po2411 = n339;
  assign po2412 = n338;
  assign po2413 = n337;
  assign po2414 = n336;
  assign po2415 = n335;
  assign po2416 = n334;
  assign po2417 = n333;
  assign po2418 = n332;
  assign po2419 = n331;
  assign po2420 = n330;
  assign po2421 = n329;
  assign po2422 = n328;
  assign po2423 = n327;
  assign po2424 = n326;
  assign po2425 = n325;
  assign po2426 = n324;
  assign po2427 = n323;
  assign po2428 = n322;
  assign po2429 = n321;
  assign po2430 = n384;
  assign po2431 = n383;
  assign po2432 = n382;
  assign po2433 = n381;
  assign po2434 = n380;
  assign po2435 = n379;
  assign po2436 = n378;
  assign po2437 = n377;
  assign po2438 = n376;
  assign po2439 = n375;
  assign po2440 = n374;
  assign po2441 = n373;
  assign po2442 = n372;
  assign po2443 = n371;
  assign po2444 = n370;
  assign po2445 = n369;
  assign po2446 = n368;
  assign po2447 = n367;
  assign po2448 = n366;
  assign po2449 = n365;
  assign po2450 = n364;
  assign po2451 = n363;
  assign po2452 = n362;
  assign po2453 = n361;
  assign po2454 = n360;
  assign po2455 = n359;
  assign po2456 = n358;
  assign po2457 = n357;
  assign po2458 = n356;
  assign po2459 = n355;
  assign po2460 = n354;
  assign po2461 = n353;
  assign po2462 = n416;
  assign po2463 = n415;
  assign po2464 = n414;
  assign po2465 = n413;
  assign po2466 = n412;
  assign po2467 = n411;
  assign po2468 = n410;
  assign po2469 = n409;
  assign po2470 = n408;
  assign po2471 = n407;
  assign po2472 = n406;
  assign po2473 = n405;
  assign po2474 = n404;
  assign po2475 = n403;
  assign po2476 = n402;
  assign po2477 = n401;
  assign po2478 = n400;
  assign po2479 = n399;
  assign po2480 = n398;
  assign po2481 = n397;
  assign po2482 = n396;
  assign po2483 = n395;
  assign po2484 = n394;
  assign po2485 = n393;
  assign po2486 = n392;
  assign po2487 = n391;
  assign po2488 = n390;
  assign po2489 = n389;
  assign po2490 = n388;
  assign po2491 = n387;
  assign po2492 = n386;
  assign po2493 = n385;
  assign po2494 = n448;
  assign po2495 = n447;
  assign po2496 = n446;
  assign po2497 = n445;
  assign po2498 = n444;
  assign po2499 = n443;
  assign po2500 = n442;
  assign po2501 = n441;
  assign po2502 = n440;
  assign po2503 = n439;
  assign po2504 = n438;
  assign po2505 = n437;
  assign po2506 = n436;
  assign po2507 = n435;
  assign po2508 = n434;
  assign po2509 = n433;
  assign po2510 = n432;
  assign po2511 = n431;
  assign po2512 = n430;
  assign po2513 = n429;
  assign po2514 = n428;
  assign po2515 = n427;
  assign po2516 = n426;
  assign po2517 = n425;
  assign po2518 = n424;
  assign po2519 = n423;
  assign po2520 = n422;
  assign po2521 = n421;
  assign po2522 = n420;
  assign po2523 = n419;
  assign po2524 = n418;
  assign po2525 = n417;
  assign po2526 = n480;
  assign po2527 = n479;
  assign po2528 = n478;
  assign po2529 = n477;
  assign po2530 = n476;
  assign po2531 = n475;
  assign po2532 = n474;
  assign po2533 = n473;
  assign po2534 = n472;
  assign po2535 = n471;
  assign po2536 = n470;
  assign po2537 = n469;
  assign po2538 = n468;
  assign po2539 = n467;
  assign po2540 = n466;
  assign po2541 = n465;
  assign po2542 = n464;
  assign po2543 = n463;
  assign po2544 = n462;
  assign po2545 = n461;
  assign po2546 = n460;
  assign po2547 = n459;
  assign po2548 = n458;
  assign po2549 = n457;
  assign po2550 = n456;
  assign po2551 = n455;
  assign po2552 = n454;
  assign po2553 = n453;
  assign po2554 = n452;
  assign po2555 = n451;
  assign po2556 = n450;
  assign po2557 = n449;
  assign po2558 = n512;
  assign po2559 = n511;
  assign po2560 = n510;
  assign po2561 = n509;
  assign po2562 = n508;
  assign po2563 = n507;
  assign po2564 = n506;
  assign po2565 = n505;
  assign po2566 = n504;
  assign po2567 = n503;
  assign po2568 = n502;
  assign po2569 = n501;
  assign po2570 = n500;
  assign po2571 = n499;
  assign po2572 = n498;
  assign po2573 = n497;
  assign po2574 = n496;
  assign po2575 = n495;
  assign po2576 = n494;
  assign po2577 = n493;
  assign po2578 = n492;
  assign po2579 = n491;
  assign po2580 = n490;
  assign po2581 = n489;
  assign po2582 = n488;
  assign po2583 = n487;
  assign po2584 = n486;
  assign po2585 = n485;
  assign po2586 = n484;
  assign po2587 = n483;
  assign po2588 = n482;
  assign po2589 = n481;
  assign po2590 = n544;
  assign po2591 = n543;
  assign po2592 = n542;
  assign po2593 = n541;
  assign po2594 = n540;
  assign po2595 = n539;
  assign po2596 = n538;
  assign po2597 = n537;
  assign po2598 = n536;
  assign po2599 = n535;
  assign po2600 = n534;
  assign po2601 = n533;
  assign po2602 = n532;
  assign po2603 = n531;
  assign po2604 = n530;
  assign po2605 = n529;
  assign po2606 = n528;
  assign po2607 = n527;
  assign po2608 = n526;
  assign po2609 = n525;
  assign po2610 = n524;
  assign po2611 = n523;
  assign po2612 = n522;
  assign po2613 = n521;
  assign po2614 = n520;
  assign po2615 = n519;
  assign po2616 = n518;
  assign po2617 = n517;
  assign po2618 = n516;
  assign po2619 = n515;
  assign po2620 = n514;
  assign po2621 = n513;
  assign po2622 = n576;
  assign po2623 = n575;
  assign po2624 = n574;
  assign po2625 = n573;
  assign po2626 = n572;
  assign po2627 = n571;
  assign po2628 = n570;
  assign po2629 = n569;
  assign po2630 = n568;
  assign po2631 = n567;
  assign po2632 = n566;
  assign po2633 = n565;
  assign po2634 = n564;
  assign po2635 = n563;
  assign po2636 = n562;
  assign po2637 = n561;
  assign po2638 = n560;
  assign po2639 = n559;
  assign po2640 = n558;
  assign po2641 = n557;
  assign po2642 = n556;
  assign po2643 = n555;
  assign po2644 = n554;
  assign po2645 = n553;
  assign po2646 = n552;
  assign po2647 = n551;
  assign po2648 = n550;
  assign po2649 = n549;
  assign po2650 = n548;
  assign po2651 = n547;
  assign po2652 = n546;
  assign po2653 = n545;
  assign po2654 = n608;
  assign po2655 = n607;
  assign po2656 = n606;
  assign po2657 = n605;
  assign po2658 = n604;
  assign po2659 = n603;
  assign po2660 = n602;
  assign po2661 = n601;
  assign po2662 = n600;
  assign po2663 = n599;
  assign po2664 = n598;
  assign po2665 = n597;
  assign po2666 = n596;
  assign po2667 = n595;
  assign po2668 = n594;
  assign po2669 = n593;
  assign po2670 = n592;
  assign po2671 = n591;
  assign po2672 = n590;
  assign po2673 = n589;
  assign po2674 = n588;
  assign po2675 = n587;
  assign po2676 = n586;
  assign po2677 = n585;
  assign po2678 = n584;
  assign po2679 = n583;
  assign po2680 = n582;
  assign po2681 = n581;
  assign po2682 = n580;
  assign po2683 = n579;
  assign po2684 = n578;
  assign po2685 = n577;
  assign po2686 = n640;
  assign po2687 = n639;
  assign po2688 = n638;
  assign po2689 = n637;
  assign po2690 = n636;
  assign po2691 = n635;
  assign po2692 = n634;
  assign po2693 = n633;
  assign po2694 = n632;
  assign po2695 = n631;
  assign po2696 = n630;
  assign po2697 = n629;
  assign po2698 = n628;
  assign po2699 = n627;
  assign po2700 = n626;
  assign po2701 = n625;
  assign po2702 = n624;
  assign po2703 = n623;
  assign po2704 = n622;
  assign po2705 = n621;
  assign po2706 = n620;
  assign po2707 = n619;
  assign po2708 = n618;
  assign po2709 = n617;
  assign po2710 = n616;
  assign po2711 = n615;
  assign po2712 = n614;
  assign po2713 = n613;
  assign po2714 = n612;
  assign po2715 = n611;
  assign po2716 = n610;
  assign po2717 = n609;
  assign po2718 = n672;
  assign po2719 = n671;
  assign po2720 = n670;
  assign po2721 = n669;
  assign po2722 = n668;
  assign po2723 = n667;
  assign po2724 = n666;
  assign po2725 = n665;
  assign po2726 = n664;
  assign po2727 = n663;
  assign po2728 = n662;
  assign po2729 = n661;
  assign po2730 = n660;
  assign po2731 = n659;
  assign po2732 = n658;
  assign po2733 = n657;
  assign po2734 = n656;
  assign po2735 = n655;
  assign po2736 = n654;
  assign po2737 = n653;
  assign po2738 = n652;
  assign po2739 = n651;
  assign po2740 = n650;
  assign po2741 = n649;
  assign po2742 = n648;
  assign po2743 = n647;
  assign po2744 = n646;
  assign po2745 = n645;
  assign po2746 = n644;
  assign po2747 = n643;
  assign po2748 = n642;
  assign po2749 = n641;
  assign po2750 = n704;
  assign po2751 = n703;
  assign po2752 = n702;
  assign po2753 = n701;
  assign po2754 = n700;
  assign po2755 = n699;
  assign po2756 = n698;
  assign po2757 = n697;
  assign po2758 = n696;
  assign po2759 = n695;
  assign po2760 = n694;
  assign po2761 = n693;
  assign po2762 = n692;
  assign po2763 = n691;
  assign po2764 = n690;
  assign po2765 = n689;
  assign po2766 = n688;
  assign po2767 = n687;
  assign po2768 = n686;
  assign po2769 = n685;
  assign po2770 = n684;
  assign po2771 = n683;
  assign po2772 = n682;
  assign po2773 = n681;
  assign po2774 = n680;
  assign po2775 = n679;
  assign po2776 = n678;
  assign po2777 = n677;
  assign po2778 = n676;
  assign po2779 = n675;
  assign po2780 = n674;
  assign po2781 = n673;
  assign po2782 = n736;
  assign po2783 = n735;
  assign po2784 = n734;
  assign po2785 = n733;
  assign po2786 = n732;
  assign po2787 = n731;
  assign po2788 = n730;
  assign po2789 = n729;
  assign po2790 = n728;
  assign po2791 = n727;
  assign po2792 = n726;
  assign po2793 = n725;
  assign po2794 = n724;
  assign po2795 = n723;
  assign po2796 = n722;
  assign po2797 = n721;
  assign po2798 = n720;
  assign po2799 = n719;
  assign po2800 = n718;
  assign po2801 = n717;
  assign po2802 = n716;
  assign po2803 = n715;
  assign po2804 = n714;
  assign po2805 = n713;
  assign po2806 = n712;
  assign po2807 = n711;
  assign po2808 = n710;
  assign po2809 = n709;
  assign po2810 = n708;
  assign po2811 = n707;
  assign po2812 = n706;
  assign po2813 = n705;
  assign po2814 = n768;
  assign po2815 = n767;
  assign po2816 = n766;
  assign po2817 = n765;
  assign po2818 = n764;
  assign po2819 = n763;
  assign po2820 = n762;
  assign po2821 = n761;
  assign po2822 = n760;
  assign po2823 = n759;
  assign po2824 = n758;
  assign po2825 = n757;
  assign po2826 = n756;
  assign po2827 = n755;
  assign po2828 = n754;
  assign po2829 = n753;
  assign po2830 = n752;
  assign po2831 = n751;
  assign po2832 = n750;
  assign po2833 = n749;
  assign po2834 = n748;
  assign po2835 = n747;
  assign po2836 = n746;
  assign po2837 = n745;
  assign po2838 = n744;
  assign po2839 = n743;
  assign po2840 = n742;
  assign po2841 = n741;
  assign po2842 = n740;
  assign po2843 = n739;
  assign po2844 = n738;
  assign po2845 = n737;
  assign po2846 = n800;
  assign po2847 = n799;
  assign po2848 = n798;
  assign po2849 = n797;
  assign po2850 = n796;
  assign po2851 = n795;
  assign po2852 = n794;
  assign po2853 = n793;
  assign po2854 = n792;
  assign po2855 = n791;
  assign po2856 = n790;
  assign po2857 = n789;
  assign po2858 = n788;
  assign po2859 = n787;
  assign po2860 = n786;
  assign po2861 = n785;
  assign po2862 = n784;
  assign po2863 = n783;
  assign po2864 = n782;
  assign po2865 = n781;
  assign po2866 = n780;
  assign po2867 = n779;
  assign po2868 = n778;
  assign po2869 = n777;
  assign po2870 = n776;
  assign po2871 = n775;
  assign po2872 = n774;
  assign po2873 = n773;
  assign po2874 = n772;
  assign po2875 = n771;
  assign po2876 = n770;
  assign po2877 = n769;
  assign po2878 = n832;
  assign po2879 = n831;
  assign po2880 = n830;
  assign po2881 = n829;
  assign po2882 = n828;
  assign po2883 = n827;
  assign po2884 = n826;
  assign po2885 = n825;
  assign po2886 = n824;
  assign po2887 = n823;
  assign po2888 = n822;
  assign po2889 = n821;
  assign po2890 = n820;
  assign po2891 = n819;
  assign po2892 = n818;
  assign po2893 = n817;
  assign po2894 = n816;
  assign po2895 = n815;
  assign po2896 = n814;
  assign po2897 = n813;
  assign po2898 = n812;
  assign po2899 = n811;
  assign po2900 = n810;
  assign po2901 = n809;
  assign po2902 = n808;
  assign po2903 = n807;
  assign po2904 = n806;
  assign po2905 = n805;
  assign po2906 = n804;
  assign po2907 = n803;
  assign po2908 = n802;
  assign po2909 = n801;
  assign po2910 = n864;
  assign po2911 = n863;
  assign po2912 = n862;
  assign po2913 = n861;
  assign po2914 = n860;
  assign po2915 = n859;
  assign po2916 = n858;
  assign po2917 = n857;
  assign po2918 = n856;
  assign po2919 = n855;
  assign po2920 = n854;
  assign po2921 = n853;
  assign po2922 = n852;
  assign po2923 = n851;
  assign po2924 = n850;
  assign po2925 = n849;
  assign po2926 = n848;
  assign po2927 = n847;
  assign po2928 = n846;
  assign po2929 = n845;
  assign po2930 = n844;
  assign po2931 = n843;
  assign po2932 = n842;
  assign po2933 = n841;
  assign po2934 = n840;
  assign po2935 = n839;
  assign po2936 = n838;
  assign po2937 = n837;
  assign po2938 = n836;
  assign po2939 = n835;
  assign po2940 = n834;
  assign po2941 = n833;
  assign po2942 = n896;
  assign po2943 = n895;
  assign po2944 = n894;
  assign po2945 = n893;
  assign po2946 = n892;
  assign po2947 = n891;
  assign po2948 = n890;
  assign po2949 = n889;
  assign po2950 = n888;
  assign po2951 = n887;
  assign po2952 = n886;
  assign po2953 = n885;
  assign po2954 = n884;
  assign po2955 = n883;
  assign po2956 = n882;
  assign po2957 = n881;
  assign po2958 = n880;
  assign po2959 = n879;
  assign po2960 = n878;
  assign po2961 = n877;
  assign po2962 = n876;
  assign po2963 = n875;
  assign po2964 = n874;
  assign po2965 = n873;
  assign po2966 = n872;
  assign po2967 = n871;
  assign po2968 = n870;
  assign po2969 = n869;
  assign po2970 = n868;
  assign po2971 = n867;
  assign po2972 = n866;
  assign po2973 = n865;
  assign po2974 = n928;
  assign po2975 = n927;
  assign po2976 = n926;
  assign po2977 = n925;
  assign po2978 = n924;
  assign po2979 = n923;
  assign po2980 = n922;
  assign po2981 = n921;
  assign po2982 = n920;
  assign po2983 = n919;
  assign po2984 = n918;
  assign po2985 = n917;
  assign po2986 = n916;
  assign po2987 = n915;
  assign po2988 = n914;
  assign po2989 = n913;
  assign po2990 = n912;
  assign po2991 = n911;
  assign po2992 = n910;
  assign po2993 = n909;
  assign po2994 = n908;
  assign po2995 = n907;
  assign po2996 = n906;
  assign po2997 = n905;
  assign po2998 = n904;
  assign po2999 = n903;
  assign po3000 = n902;
  assign po3001 = n901;
  assign po3002 = n900;
  assign po3003 = n899;
  assign po3004 = n898;
  assign po3005 = n897;
  assign po3006 = n960;
  assign po3007 = n959;
  assign po3008 = n958;
  assign po3009 = n957;
  assign po3010 = n956;
  assign po3011 = n955;
  assign po3012 = n954;
  assign po3013 = n953;
  assign po3014 = n952;
  assign po3015 = n951;
  assign po3016 = n950;
  assign po3017 = n949;
  assign po3018 = n948;
  assign po3019 = n947;
  assign po3020 = n946;
  assign po3021 = n945;
  assign po3022 = n944;
  assign po3023 = n943;
  assign po3024 = n942;
  assign po3025 = n941;
  assign po3026 = n940;
  assign po3027 = n939;
  assign po3028 = n938;
  assign po3029 = n937;
  assign po3030 = n936;
  assign po3031 = n935;
  assign po3032 = n934;
  assign po3033 = n933;
  assign po3034 = n932;
  assign po3035 = n931;
  assign po3036 = n930;
  assign po3037 = n929;
  assign po3038 = n992;
  assign po3039 = n991;
  assign po3040 = n990;
  assign po3041 = n989;
  assign po3042 = n988;
  assign po3043 = n987;
  assign po3044 = n986;
  assign po3045 = n985;
  assign po3046 = n984;
  assign po3047 = n983;
  assign po3048 = n982;
  assign po3049 = n981;
  assign po3050 = n980;
  assign po3051 = n979;
  assign po3052 = n978;
  assign po3053 = n977;
  assign po3054 = n976;
  assign po3055 = n975;
  assign po3056 = n974;
  assign po3057 = n973;
  assign po3058 = n972;
  assign po3059 = n971;
  assign po3060 = n970;
  assign po3061 = n969;
  assign po3062 = n968;
  assign po3063 = n967;
  assign po3064 = n966;
  assign po3065 = n965;
  assign po3066 = n964;
  assign po3067 = n963;
  assign po3068 = n962;
  assign po3069 = n961;
  assign po3070 = n1024;
  assign po3071 = n1023;
  assign po3072 = n1022;
  assign po3073 = n1021;
  assign po3074 = n1020;
  assign po3075 = n1019;
  assign po3076 = n1018;
  assign po3077 = n1017;
  assign po3078 = n1016;
  assign po3079 = n1015;
  assign po3080 = n1014;
  assign po3081 = n1013;
  assign po3082 = n1012;
  assign po3083 = n1011;
  assign po3084 = n1010;
  assign po3085 = n1009;
  assign po3086 = n1008;
  assign po3087 = n1007;
  assign po3088 = n1006;
  assign po3089 = n1005;
  assign po3090 = n1004;
  assign po3091 = n1003;
  assign po3092 = n1002;
  assign po3093 = n1001;
  assign po3094 = n1000;
  assign po3095 = n999;
  assign po3096 = n998;
  assign po3097 = n997;
  assign po3098 = n996;
  assign po3099 = n995;
  assign po3100 = n994;
  assign po3101 = n993;
  assign po3102 = n1056;
  assign po3103 = n1055;
  assign po3104 = n1054;
  assign po3105 = n1053;
  assign po3106 = n1052;
  assign po3107 = n1051;
  assign po3108 = n1050;
  assign po3109 = n1049;
  assign po3110 = n1048;
  assign po3111 = n1047;
  assign po3112 = n1046;
  assign po3113 = n1045;
  assign po3114 = n1044;
  assign po3115 = n1043;
  assign po3116 = n1042;
  assign po3117 = n1041;
  assign po3118 = n1040;
  assign po3119 = n1039;
  assign po3120 = n1038;
  assign po3121 = n1037;
  assign po3122 = n1036;
  assign po3123 = n1035;
  assign po3124 = n1034;
  assign po3125 = n1033;
  assign po3126 = n1032;
  assign po3127 = n1031;
  assign po3128 = n1030;
  assign po3129 = n1029;
  assign po3130 = n1028;
  assign po3131 = n1027;
  assign po3132 = n1026;
  assign po3133 = n1025;
  assign po3134 = n1088;
  assign po3135 = n1087;
  assign po3136 = n1086;
  assign po3137 = n1085;
  assign po3138 = n1084;
  assign po3139 = n1083;
  assign po3140 = n1082;
  assign po3141 = n1081;
  assign po3142 = n1080;
  assign po3143 = n1079;
  assign po3144 = n1078;
  assign po3145 = n1077;
  assign po3146 = n1076;
  assign po3147 = n1075;
  assign po3148 = n1074;
  assign po3149 = n1073;
  assign po3150 = n1072;
  assign po3151 = n1071;
  assign po3152 = n1070;
  assign po3153 = n1069;
  assign po3154 = n1068;
  assign po3155 = n1067;
  assign po3156 = n1066;
  assign po3157 = n1065;
  assign po3158 = n1064;
  assign po3159 = n1063;
  assign po3160 = n1062;
  assign po3161 = n1061;
  assign po3162 = n1060;
  assign po3163 = n1059;
  assign po3164 = n1058;
  assign po3165 = n1057;
  assign po3166 = n1120;
  assign po3167 = n1119;
  assign po3168 = n1118;
  assign po3169 = n1117;
  assign po3170 = n1116;
  assign po3171 = n1115;
  assign po3172 = n1114;
  assign po3173 = n1113;
  assign po3174 = n1112;
  assign po3175 = n1111;
  assign po3176 = n1110;
  assign po3177 = n1109;
  assign po3178 = n1108;
  assign po3179 = n1107;
  assign po3180 = n1106;
  assign po3181 = n1105;
  assign po3182 = n1104;
  assign po3183 = n1103;
  assign po3184 = n1102;
  assign po3185 = n1101;
  assign po3186 = n1100;
  assign po3187 = n1099;
  assign po3188 = n1098;
  assign po3189 = n1097;
  assign po3190 = n1096;
  assign po3191 = n1095;
  assign po3192 = n1094;
  assign po3193 = n1093;
  assign po3194 = n1092;
  assign po3195 = n1091;
  assign po3196 = n1090;
  assign po3197 = n1089;
  assign po3198 = n1152;
  assign po3199 = n1151;
  assign po3200 = n1150;
  assign po3201 = n1149;
  assign po3202 = n1148;
  assign po3203 = n1147;
  assign po3204 = n1146;
  assign po3205 = n1145;
  assign po3206 = n1144;
  assign po3207 = n1143;
  assign po3208 = n1142;
  assign po3209 = n1141;
  assign po3210 = n1140;
  assign po3211 = n1139;
  assign po3212 = n1138;
  assign po3213 = n1137;
  assign po3214 = n1136;
  assign po3215 = n1135;
  assign po3216 = n1134;
  assign po3217 = n1133;
  assign po3218 = n1132;
  assign po3219 = n1131;
  assign po3220 = n1130;
  assign po3221 = n1129;
  assign po3222 = n1128;
  assign po3223 = n1127;
  assign po3224 = n1126;
  assign po3225 = n1125;
  assign po3226 = n1124;
  assign po3227 = n1123;
  assign po3228 = n1122;
  assign po3229 = n1121;
  assign po3230 = n1184;
  assign po3231 = n1183;
  assign po3232 = n1182;
  assign po3233 = n1181;
  assign po3234 = n1180;
  assign po3235 = n1179;
  assign po3236 = n1178;
  assign po3237 = n1177;
  assign po3238 = n1176;
  assign po3239 = n1175;
  assign po3240 = n1174;
  assign po3241 = n1173;
  assign po3242 = n1172;
  assign po3243 = n1171;
  assign po3244 = n1170;
  assign po3245 = n1169;
  assign po3246 = n1168;
  assign po3247 = n1167;
  assign po3248 = n1166;
  assign po3249 = n1165;
  assign po3250 = n1164;
  assign po3251 = n1163;
  assign po3252 = n1162;
  assign po3253 = n1161;
  assign po3254 = n1160;
  assign po3255 = n1159;
  assign po3256 = n1158;
  assign po3257 = n1157;
  assign po3258 = n1156;
  assign po3259 = n1155;
  assign po3260 = n1154;
  assign po3261 = n1153;
  assign po3262 = n1216;
  assign po3263 = n1215;
  assign po3264 = n1214;
  assign po3265 = n1213;
  assign po3266 = n1212;
  assign po3267 = n1211;
  assign po3268 = n1210;
  assign po3269 = n1209;
  assign po3270 = n1208;
  assign po3271 = n1207;
  assign po3272 = n1206;
  assign po3273 = n1205;
  assign po3274 = n1204;
  assign po3275 = n1203;
  assign po3276 = n1202;
  assign po3277 = n1201;
  assign po3278 = n1200;
  assign po3279 = n1199;
  assign po3280 = n1198;
  assign po3281 = n1197;
  assign po3282 = n1196;
  assign po3283 = n1195;
  assign po3284 = n1194;
  assign po3285 = n1193;
  assign po3286 = n1192;
  assign po3287 = n1191;
  assign po3288 = n1190;
  assign po3289 = n1189;
  assign po3290 = n1188;
  assign po3291 = n1187;
  assign po3292 = n1186;
  assign po3293 = n1185;
  assign po3294 = n1248;
  assign po3295 = n1247;
  assign po3296 = n1246;
  assign po3297 = n1245;
  assign po3298 = n1244;
  assign po3299 = n1243;
  assign po3300 = n1242;
  assign po3301 = n1241;
  assign po3302 = n1240;
  assign po3303 = n1239;
  assign po3304 = n1238;
  assign po3305 = n1237;
  assign po3306 = n1236;
  assign po3307 = n1235;
  assign po3308 = n1234;
  assign po3309 = n1233;
  assign po3310 = n1232;
  assign po3311 = n1231;
  assign po3312 = n1230;
  assign po3313 = n1229;
  assign po3314 = n1228;
  assign po3315 = n1227;
  assign po3316 = n1226;
  assign po3317 = n1225;
  assign po3318 = n1224;
  assign po3319 = n1223;
  assign po3320 = n1222;
  assign po3321 = n1221;
  assign po3322 = n1220;
  assign po3323 = n1219;
  assign po3324 = n1218;
  assign po3325 = n1217;
  assign po3326 = n1280;
  assign po3327 = n1279;
  assign po3328 = n1278;
  assign po3329 = n1277;
  assign po3330 = n1276;
  assign po3331 = n1275;
  assign po3332 = n1274;
  assign po3333 = n1273;
  assign po3334 = n1272;
  assign po3335 = n1271;
  assign po3336 = n1270;
  assign po3337 = n1269;
  assign po3338 = n1268;
  assign po3339 = n1267;
  assign po3340 = n1266;
  assign po3341 = n1265;
  assign po3342 = n1264;
  assign po3343 = n1263;
  assign po3344 = n1262;
  assign po3345 = n1261;
  assign po3346 = n1260;
  assign po3347 = n1259;
  assign po3348 = n1258;
  assign po3349 = n1257;
  assign po3350 = n1256;
  assign po3351 = n1255;
  assign po3352 = n1254;
  assign po3353 = n1253;
  assign po3354 = n1252;
  assign po3355 = n1251;
  assign po3356 = n1250;
  assign po3357 = n1249;
  assign po3358 = n1312;
  assign po3359 = n1311;
  assign po3360 = n1310;
  assign po3361 = n1309;
  assign po3362 = n1308;
  assign po3363 = n1307;
  assign po3364 = n1306;
  assign po3365 = n1305;
  assign po3366 = n1304;
  assign po3367 = n1303;
  assign po3368 = n1302;
  assign po3369 = n1301;
  assign po3370 = n1300;
  assign po3371 = n1299;
  assign po3372 = n1298;
  assign po3373 = n1297;
  assign po3374 = n1296;
  assign po3375 = n1295;
  assign po3376 = n1294;
  assign po3377 = n1293;
  assign po3378 = n1292;
  assign po3379 = n1291;
  assign po3380 = n1290;
  assign po3381 = n1289;
  assign po3382 = n1288;
  assign po3383 = n1287;
  assign po3384 = n1286;
  assign po3385 = n1285;
  assign po3386 = n1284;
  assign po3387 = n1283;
  assign po3388 = n1282;
  assign po3389 = n1281;
  assign po3390 = n1344;
  assign po3391 = n1343;
  assign po3392 = n1342;
  assign po3393 = n1341;
  assign po3394 = n1340;
  assign po3395 = n1339;
  assign po3396 = n1338;
  assign po3397 = n1337;
  assign po3398 = n1336;
  assign po3399 = n1335;
  assign po3400 = n1334;
  assign po3401 = n1333;
  assign po3402 = n1332;
  assign po3403 = n1331;
  assign po3404 = n1330;
  assign po3405 = n1329;
  assign po3406 = n1328;
  assign po3407 = n1327;
  assign po3408 = n1326;
  assign po3409 = n1325;
  assign po3410 = n1324;
  assign po3411 = n1323;
  assign po3412 = n1322;
  assign po3413 = n1321;
  assign po3414 = n1320;
  assign po3415 = n1319;
  assign po3416 = n1318;
  assign po3417 = n1317;
  assign po3418 = n1316;
  assign po3419 = n1315;
  assign po3420 = n1314;
  assign po3421 = n1313;
  assign po3422 = n1376;
  assign po3423 = n1375;
  assign po3424 = n1374;
  assign po3425 = n1373;
  assign po3426 = n1372;
  assign po3427 = n1371;
  assign po3428 = n1370;
  assign po3429 = n1369;
  assign po3430 = n1368;
  assign po3431 = n1367;
  assign po3432 = n1366;
  assign po3433 = n1365;
  assign po3434 = n1364;
  assign po3435 = n1363;
  assign po3436 = n1362;
  assign po3437 = n1361;
  assign po3438 = n1360;
  assign po3439 = n1359;
  assign po3440 = n1358;
  assign po3441 = n1357;
  assign po3442 = n1356;
  assign po3443 = n1355;
  assign po3444 = n1354;
  assign po3445 = n1353;
  assign po3446 = n1352;
  assign po3447 = n1351;
  assign po3448 = n1350;
  assign po3449 = n1349;
  assign po3450 = n1348;
  assign po3451 = n1347;
  assign po3452 = n1346;
  assign po3453 = n1345;
  assign po3454 = n1408;
  assign po3455 = n1407;
  assign po3456 = n1406;
  assign po3457 = n1405;
  assign po3458 = n1404;
  assign po3459 = n1403;
  assign po3460 = n1402;
  assign po3461 = n1401;
  assign po3462 = n1400;
  assign po3463 = n1399;
  assign po3464 = n1398;
  assign po3465 = n1397;
  assign po3466 = n1396;
  assign po3467 = n1395;
  assign po3468 = n1394;
  assign po3469 = n1393;
  assign po3470 = n1392;
  assign po3471 = n1391;
  assign po3472 = n1390;
  assign po3473 = n1389;
  assign po3474 = n1388;
  assign po3475 = n1387;
  assign po3476 = n1386;
  assign po3477 = n1385;
  assign po3478 = n1384;
  assign po3479 = n1383;
  assign po3480 = n1382;
  assign po3481 = n1381;
  assign po3482 = n1380;
  assign po3483 = n1379;
  assign po3484 = n1378;
  assign po3485 = n1377;
  assign po3486 = n1440;
  assign po3487 = n1439;
  assign po3488 = n1438;
  assign po3489 = n1437;
  assign po3490 = n1436;
  assign po3491 = n1435;
  assign po3492 = n1434;
  assign po3493 = n1433;
  assign po3494 = n1432;
  assign po3495 = n1431;
  assign po3496 = n1430;
  assign po3497 = n1429;
  assign po3498 = n1428;
  assign po3499 = n1427;
  assign po3500 = n1426;
  assign po3501 = n1425;
  assign po3502 = n1424;
  assign po3503 = n1423;
  assign po3504 = n1422;
  assign po3505 = n1421;
  assign po3506 = n1420;
  assign po3507 = n1419;
  assign po3508 = n1418;
  assign po3509 = n1417;
  assign po3510 = n1416;
  assign po3511 = n1415;
  assign po3512 = n1414;
  assign po3513 = n1413;
  assign po3514 = n1412;
  assign po3515 = n1411;
  assign po3516 = n1410;
  assign po3517 = n1409;
  assign po3518 = n1472;
  assign po3519 = n1471;
  assign po3520 = n1470;
  assign po3521 = n1469;
  assign po3522 = n1468;
  assign po3523 = n1467;
  assign po3524 = n1466;
  assign po3525 = n1465;
  assign po3526 = n1464;
  assign po3527 = n1463;
  assign po3528 = n1462;
  assign po3529 = n1461;
  assign po3530 = n1460;
  assign po3531 = n1459;
  assign po3532 = n1458;
  assign po3533 = n1457;
  assign po3534 = n1456;
  assign po3535 = n1455;
  assign po3536 = n1454;
  assign po3537 = n1453;
  assign po3538 = n1452;
  assign po3539 = n1451;
  assign po3540 = n1450;
  assign po3541 = n1449;
  assign po3542 = n1448;
  assign po3543 = n1447;
  assign po3544 = n1446;
  assign po3545 = n1445;
  assign po3546 = n1444;
  assign po3547 = n1443;
  assign po3548 = n1442;
  assign po3549 = n1441;
  assign po3550 = n1504;
  assign po3551 = n1503;
  assign po3552 = n1502;
  assign po3553 = n1501;
  assign po3554 = n1500;
  assign po3555 = n1499;
  assign po3556 = n1498;
  assign po3557 = n1497;
  assign po3558 = n1496;
  assign po3559 = n1495;
  assign po3560 = n1494;
  assign po3561 = n1493;
  assign po3562 = n1492;
  assign po3563 = n1491;
  assign po3564 = n1490;
  assign po3565 = n1489;
  assign po3566 = n1488;
  assign po3567 = n1487;
  assign po3568 = n1486;
  assign po3569 = n1485;
  assign po3570 = n1484;
  assign po3571 = n1483;
  assign po3572 = n1482;
  assign po3573 = n1481;
  assign po3574 = n1480;
  assign po3575 = n1479;
  assign po3576 = n1478;
  assign po3577 = n1477;
  assign po3578 = n1476;
  assign po3579 = n1475;
  assign po3580 = n1474;
  assign po3581 = n1473;
  assign po3582 = n1536;
  assign po3583 = n1535;
  assign po3584 = n1534;
  assign po3585 = n1533;
  assign po3586 = n1532;
  assign po3587 = n1531;
  assign po3588 = n1530;
  assign po3589 = n1529;
  assign po3590 = n1528;
  assign po3591 = n1527;
  assign po3592 = n1526;
  assign po3593 = n1525;
  assign po3594 = n1524;
  assign po3595 = n1523;
  assign po3596 = n1522;
  assign po3597 = n1521;
  assign po3598 = n1520;
  assign po3599 = n1519;
  assign po3600 = n1518;
  assign po3601 = n1517;
  assign po3602 = n1516;
  assign po3603 = n1515;
  assign po3604 = n1514;
  assign po3605 = n1513;
  assign po3606 = n1512;
  assign po3607 = n1511;
  assign po3608 = n1510;
  assign po3609 = n1509;
  assign po3610 = n1508;
  assign po3611 = n1507;
  assign po3612 = n1506;
  assign po3613 = n1505;
  assign po3614 = n1568;
  assign po3615 = n1567;
  assign po3616 = n1566;
  assign po3617 = n1565;
  assign po3618 = n1564;
  assign po3619 = n1563;
  assign po3620 = n1562;
  assign po3621 = n1561;
  assign po3622 = n1560;
  assign po3623 = n1559;
  assign po3624 = n1558;
  assign po3625 = n1557;
  assign po3626 = n1556;
  assign po3627 = n1555;
  assign po3628 = n1554;
  assign po3629 = n1553;
  assign po3630 = n1552;
  assign po3631 = n1551;
  assign po3632 = n1550;
  assign po3633 = n1549;
  assign po3634 = n1548;
  assign po3635 = n1547;
  assign po3636 = n1546;
  assign po3637 = n1545;
  assign po3638 = n1544;
  assign po3639 = n1543;
  assign po3640 = n1542;
  assign po3641 = n1541;
  assign po3642 = n1540;
  assign po3643 = n1539;
  assign po3644 = n1538;
  assign po3645 = n1537;
  assign po3646 = n1600;
  assign po3647 = n1599;
  assign po3648 = n1598;
  assign po3649 = n1597;
  assign po3650 = n1596;
  assign po3651 = n1595;
  assign po3652 = n1594;
  assign po3653 = n1593;
  assign po3654 = n1592;
  assign po3655 = n1591;
  assign po3656 = n1590;
  assign po3657 = n1589;
  assign po3658 = n1588;
  assign po3659 = n1587;
  assign po3660 = n1586;
  assign po3661 = n1585;
  assign po3662 = n1584;
  assign po3663 = n1583;
  assign po3664 = n1582;
  assign po3665 = n1581;
  assign po3666 = n1580;
  assign po3667 = n1579;
  assign po3668 = n1578;
  assign po3669 = n1577;
  assign po3670 = n1576;
  assign po3671 = n1575;
  assign po3672 = n1574;
  assign po3673 = n1573;
  assign po3674 = n1572;
  assign po3675 = n1571;
  assign po3676 = n1570;
  assign po3677 = n1569;
  assign po3678 = n1632;
  assign po3679 = n1631;
  assign po3680 = n1630;
  assign po3681 = n1629;
  assign po3682 = n1628;
  assign po3683 = n1627;
  assign po3684 = n1626;
  assign po3685 = n1625;
  assign po3686 = n1624;
  assign po3687 = n1623;
  assign po3688 = n1622;
  assign po3689 = n1621;
  assign po3690 = n1620;
  assign po3691 = n1619;
  assign po3692 = n1618;
  assign po3693 = n1617;
  assign po3694 = n1616;
  assign po3695 = n1615;
  assign po3696 = n1614;
  assign po3697 = n1613;
  assign po3698 = n1612;
  assign po3699 = n1611;
  assign po3700 = n1610;
  assign po3701 = n1609;
  assign po3702 = n1608;
  assign po3703 = n1607;
  assign po3704 = n1606;
  assign po3705 = n1605;
  assign po3706 = n1604;
  assign po3707 = n1603;
  assign po3708 = n1602;
  assign po3709 = n1601;
  assign po3710 = n1664;
  assign po3711 = n1663;
  assign po3712 = n1662;
  assign po3713 = n1661;
  assign po3714 = n1660;
  assign po3715 = n1659;
  assign po3716 = n1658;
  assign po3717 = n1657;
  assign po3718 = n1656;
  assign po3719 = n1655;
  assign po3720 = n1654;
  assign po3721 = n1653;
  assign po3722 = n1652;
  assign po3723 = n1651;
  assign po3724 = n1650;
  assign po3725 = n1649;
  assign po3726 = n1648;
  assign po3727 = n1647;
  assign po3728 = n1646;
  assign po3729 = n1645;
  assign po3730 = n1644;
  assign po3731 = n1643;
  assign po3732 = n1642;
  assign po3733 = n1641;
  assign po3734 = n1640;
  assign po3735 = n1639;
  assign po3736 = n1638;
  assign po3737 = n1637;
  assign po3738 = n1636;
  assign po3739 = n1635;
  assign po3740 = n1634;
  assign po3741 = n1633;
  assign po3742 = n1696;
  assign po3743 = n1695;
  assign po3744 = n1694;
  assign po3745 = n1693;
  assign po3746 = n1692;
  assign po3747 = n1691;
  assign po3748 = n1690;
  assign po3749 = n1689;
  assign po3750 = n1688;
  assign po3751 = n1687;
  assign po3752 = n1686;
  assign po3753 = n1685;
  assign po3754 = n1684;
  assign po3755 = n1683;
  assign po3756 = n1682;
  assign po3757 = n1681;
  assign po3758 = n1680;
  assign po3759 = n1679;
  assign po3760 = n1678;
  assign po3761 = n1677;
  assign po3762 = n1676;
  assign po3763 = n1675;
  assign po3764 = n1674;
  assign po3765 = n1673;
  assign po3766 = n1672;
  assign po3767 = n1671;
  assign po3768 = n1670;
  assign po3769 = n1669;
  assign po3770 = n1668;
  assign po3771 = n1667;
  assign po3772 = n1666;
  assign po3773 = n1665;
  assign po3774 = n1728;
  assign po3775 = n1727;
  assign po3776 = n1726;
  assign po3777 = n1725;
  assign po3778 = n1724;
  assign po3779 = n1723;
  assign po3780 = n1722;
  assign po3781 = n1721;
  assign po3782 = n1720;
  assign po3783 = n1719;
  assign po3784 = n1718;
  assign po3785 = n1717;
  assign po3786 = n1716;
  assign po3787 = n1715;
  assign po3788 = n1714;
  assign po3789 = n1713;
  assign po3790 = n1712;
  assign po3791 = n1711;
  assign po3792 = n1710;
  assign po3793 = n1709;
  assign po3794 = n1708;
  assign po3795 = n1707;
  assign po3796 = n1706;
  assign po3797 = n1705;
  assign po3798 = n1704;
  assign po3799 = n1703;
  assign po3800 = n1702;
  assign po3801 = n1701;
  assign po3802 = n1700;
  assign po3803 = n1699;
  assign po3804 = n1698;
  assign po3805 = n1697;
  assign po3806 = n1760;
  assign po3807 = n1759;
  assign po3808 = n1758;
  assign po3809 = n1757;
  assign po3810 = n1756;
  assign po3811 = n1755;
  assign po3812 = n1754;
  assign po3813 = n1753;
  assign po3814 = n1752;
  assign po3815 = n1751;
  assign po3816 = n1750;
  assign po3817 = n1749;
  assign po3818 = n1748;
  assign po3819 = n1747;
  assign po3820 = n1746;
  assign po3821 = n1745;
  assign po3822 = n1744;
  assign po3823 = n1743;
  assign po3824 = n1742;
  assign po3825 = n1741;
  assign po3826 = n1740;
  assign po3827 = n1739;
  assign po3828 = n1738;
  assign po3829 = n1737;
  assign po3830 = n1736;
  assign po3831 = n1735;
  assign po3832 = n1734;
  assign po3833 = n1733;
  assign po3834 = n1732;
  assign po3835 = n1731;
  assign po3836 = n1730;
  assign po3837 = n1729;
  assign po3838 = n1792;
  assign po3839 = n1791;
  assign po3840 = n1790;
  assign po3841 = n1789;
  assign po3842 = n1788;
  assign po3843 = n1787;
  assign po3844 = n1786;
  assign po3845 = n1785;
  assign po3846 = n1784;
  assign po3847 = n1783;
  assign po3848 = n1782;
  assign po3849 = n1781;
  assign po3850 = n1780;
  assign po3851 = n1779;
  assign po3852 = n1778;
  assign po3853 = n1777;
  assign po3854 = n1776;
  assign po3855 = n1775;
  assign po3856 = n1774;
  assign po3857 = n1773;
  assign po3858 = n1772;
  assign po3859 = n1771;
  assign po3860 = n1770;
  assign po3861 = n1769;
  assign po3862 = n1768;
  assign po3863 = n1767;
  assign po3864 = n1766;
  assign po3865 = n1765;
  assign po3866 = n1764;
  assign po3867 = n1763;
  assign po3868 = n1762;
  assign po3869 = n1761;
  assign po3870 = n1824;
  assign po3871 = n1823;
  assign po3872 = n1822;
  assign po3873 = n1821;
  assign po3874 = n1820;
  assign po3875 = n1819;
  assign po3876 = n1818;
  assign po3877 = n1817;
  assign po3878 = n1816;
  assign po3879 = n1815;
  assign po3880 = n1814;
  assign po3881 = n1813;
  assign po3882 = n1812;
  assign po3883 = n1811;
  assign po3884 = n1810;
  assign po3885 = n1809;
  assign po3886 = n1808;
  assign po3887 = n1807;
  assign po3888 = n1806;
  assign po3889 = n1805;
  assign po3890 = n1804;
  assign po3891 = n1803;
  assign po3892 = n1802;
  assign po3893 = n1801;
  assign po3894 = n1800;
  assign po3895 = n1799;
  assign po3896 = n1798;
  assign po3897 = n1797;
  assign po3898 = n1796;
  assign po3899 = n1795;
  assign po3900 = n1794;
  assign po3901 = n1793;
  assign po3902 = n1856;
  assign po3903 = n1855;
  assign po3904 = n1854;
  assign po3905 = n1853;
  assign po3906 = n1852;
  assign po3907 = n1851;
  assign po3908 = n1850;
  assign po3909 = n1849;
  assign po3910 = n1848;
  assign po3911 = n1847;
  assign po3912 = n1846;
  assign po3913 = n1845;
  assign po3914 = n1844;
  assign po3915 = n1843;
  assign po3916 = n1842;
  assign po3917 = n1841;
  assign po3918 = n1840;
  assign po3919 = n1839;
  assign po3920 = n1838;
  assign po3921 = n1837;
  assign po3922 = n1836;
  assign po3923 = n1835;
  assign po3924 = n1834;
  assign po3925 = n1833;
  assign po3926 = n1832;
  assign po3927 = n1831;
  assign po3928 = n1830;
  assign po3929 = n1829;
  assign po3930 = n1828;
  assign po3931 = n1827;
  assign po3932 = n1826;
  assign po3933 = n1825;
  assign po3934 = n1888;
  assign po3935 = n1887;
  assign po3936 = n1886;
  assign po3937 = n1885;
  assign po3938 = n1884;
  assign po3939 = n1883;
  assign po3940 = n1882;
  assign po3941 = n1881;
  assign po3942 = n1880;
  assign po3943 = n1879;
  assign po3944 = n1878;
  assign po3945 = n1877;
  assign po3946 = n1876;
  assign po3947 = n1875;
  assign po3948 = n1874;
  assign po3949 = n1873;
  assign po3950 = n1872;
  assign po3951 = n1871;
  assign po3952 = n1870;
  assign po3953 = n1869;
  assign po3954 = n1868;
  assign po3955 = n1867;
  assign po3956 = n1866;
  assign po3957 = n1865;
  assign po3958 = n1864;
  assign po3959 = n1863;
  assign po3960 = n1862;
  assign po3961 = n1861;
  assign po3962 = n1860;
  assign po3963 = n1859;
  assign po3964 = n1858;
  assign po3965 = n1857;
  assign po3966 = n1920;
  assign po3967 = n1919;
  assign po3968 = n1918;
  assign po3969 = n1917;
  assign po3970 = n1916;
  assign po3971 = n1915;
  assign po3972 = n1914;
  assign po3973 = n1913;
  assign po3974 = n1912;
  assign po3975 = n1911;
  assign po3976 = n1910;
  assign po3977 = n1909;
  assign po3978 = n1908;
  assign po3979 = n1907;
  assign po3980 = n1906;
  assign po3981 = n1905;
  assign po3982 = n1904;
  assign po3983 = n1903;
  assign po3984 = n1902;
  assign po3985 = n1901;
  assign po3986 = n1900;
  assign po3987 = n1899;
  assign po3988 = n1898;
  assign po3989 = n1897;
  assign po3990 = n1896;
  assign po3991 = n1895;
  assign po3992 = n1894;
  assign po3993 = n1893;
  assign po3994 = n1892;
  assign po3995 = n1891;
  assign po3996 = n1890;
  assign po3997 = n1889;
  assign po3998 = n1952;
  assign po3999 = n1951;
  assign po4000 = n1950;
  assign po4001 = n1949;
  assign po4002 = n1948;
  assign po4003 = n1947;
  assign po4004 = n1946;
  assign po4005 = n1945;
  assign po4006 = n1944;
  assign po4007 = n1943;
  assign po4008 = n1942;
  assign po4009 = n1941;
  assign po4010 = n1940;
  assign po4011 = n1939;
  assign po4012 = n1938;
  assign po4013 = n1937;
  assign po4014 = n1936;
  assign po4015 = n1935;
  assign po4016 = n1934;
  assign po4017 = n1933;
  assign po4018 = n1932;
  assign po4019 = n1931;
  assign po4020 = n1930;
  assign po4021 = n1929;
  assign po4022 = n1928;
  assign po4023 = n1927;
  assign po4024 = n1926;
  assign po4025 = n1925;
  assign po4026 = n1924;
  assign po4027 = n1923;
  assign po4028 = n1922;
  assign po4029 = n1921;
  assign po4030 = n1984;
  assign po4031 = n1983;
  assign po4032 = n1982;
  assign po4033 = n1981;
  assign po4034 = n1980;
  assign po4035 = n1979;
  assign po4036 = n1978;
  assign po4037 = n1977;
  assign po4038 = n1976;
  assign po4039 = n1975;
  assign po4040 = n1974;
  assign po4041 = n1973;
  assign po4042 = n1972;
  assign po4043 = n1971;
  assign po4044 = n1970;
  assign po4045 = n1969;
  assign po4046 = n1968;
  assign po4047 = n1967;
  assign po4048 = n1966;
  assign po4049 = n1965;
  assign po4050 = n1964;
  assign po4051 = n1963;
  assign po4052 = n1962;
  assign po4053 = n1961;
  assign po4054 = n1960;
  assign po4055 = n1959;
  assign po4056 = n1958;
  assign po4057 = n1957;
  assign po4058 = n1956;
  assign po4059 = n1955;
  assign po4060 = n1954;
  assign po4061 = n1953;
  assign po4062 = n2016;
  assign po4063 = n2015;
  assign po4064 = n2014;
  assign po4065 = n2013;
  assign po4066 = n2012;
  assign po4067 = n2011;
  assign po4068 = n2010;
  assign po4069 = n2009;
  assign po4070 = n2008;
  assign po4071 = n2007;
  assign po4072 = n2006;
  assign po4073 = n2005;
  assign po4074 = n2004;
  assign po4075 = n2003;
  assign po4076 = n2002;
  assign po4077 = n2001;
  assign po4078 = n2000;
  assign po4079 = n1999;
  assign po4080 = n1998;
  assign po4081 = n1997;
  assign po4082 = n1996;
  assign po4083 = n1995;
  assign po4084 = n1994;
  assign po4085 = n1993;
  assign po4086 = n1992;
  assign po4087 = n1991;
  assign po4088 = n1990;
  assign po4089 = n1989;
  assign po4090 = n1988;
  assign po4091 = n1987;
  assign po4092 = n1986;
  assign po4093 = n1985;
  assign po4094 = n2048;
  assign po4095 = n2047;
  assign po4096 = n2046;
  assign po4097 = n2045;
  assign po4098 = n2044;
  assign po4099 = n2043;
  assign po4100 = n2042;
  assign po4101 = n2041;
  assign po4102 = n2040;
  assign po4103 = n2039;
  assign po4104 = n2038;
  assign po4105 = n2037;
  assign po4106 = n2036;
  assign po4107 = n2035;
  assign po4108 = n2034;
  assign po4109 = n2033;
  assign po4110 = n2032;
  assign po4111 = n2031;
  assign po4112 = n2030;
  assign po4113 = n2029;
  assign po4114 = n2028;
  assign po4115 = n2027;
  assign po4116 = n2026;
  assign po4117 = n2025;
  assign po4118 = n2024;
  assign po4119 = n2023;
  assign po4120 = n2022;
  assign po4121 = n2021;
  assign po4122 = n2020;
  assign po4123 = n2019;
  assign po4124 = n2018;
  assign po4125 = n2017;
  assign po4126 = new_n5441;
  assign po4127 = new_n5442;
  assign po4128 = new_n5443;
  assign po4129 = new_n5444;
  assign po4130 = new_n5445;
  assign po4131 = new_n5446;
  assign po4132 = new_n5447;
  assign po4133 = new_n5448;
  assign po4134 = new_n5452;
  assign po4135 = new_n5453;
  assign po4136 = new_n5454;
  assign po4137 = new_n5455;
  assign po4138 = new_n5456;
  assign po4139 = new_n5457;
  assign po4140 = new_n5458;
  assign po4141 = new_n5459;
  assign po4142 = new_n5465;
  assign po4143 = new_n5466;
  assign po4144 = new_n5467;
  assign po4145 = new_n5468;
  assign po4146 = new_n5469;
  assign po4147 = new_n5470;
  assign po4148 = new_n5471;
  assign po4149 = new_n5472;
  assign po4150 = new_n5475;
  assign po4151 = new_n5476;
  assign po4152 = new_n5477;
  assign po4153 = new_n5478;
  assign po4154 = new_n5479;
  assign po4155 = new_n5480;
  assign po4156 = new_n5481;
  assign po4157 = new_n5482;
  assign po4158 = new_n5492;
  assign po4159 = new_n5493;
  assign po4160 = new_n5494;
  assign po4161 = new_n5495;
  assign po4162 = new_n5496;
  assign po4163 = new_n5497;
  assign po4164 = new_n5498;
  assign po4165 = new_n5499;
  assign po4166 = new_n5503;
  assign po4167 = new_n5504;
  assign po4168 = new_n5505;
  assign po4169 = new_n5506;
  assign po4170 = new_n5507;
  assign po4171 = new_n5508;
  assign po4172 = new_n5509;
  assign po4173 = new_n5510;
  assign po4174 = new_n5516;
  assign po4175 = new_n5517;
  assign po4176 = new_n5518;
  assign po4177 = new_n5519;
  assign po4178 = new_n5520;
  assign po4179 = new_n5521;
  assign po4180 = new_n5522;
  assign po4181 = new_n5523;
  assign po4182 = new_n5527;
  assign po4183 = new_n5528;
  assign po4184 = new_n5529;
  assign po4185 = new_n5530;
  assign po4186 = new_n5531;
  assign po4187 = new_n5532;
  assign po4188 = new_n5533;
  assign po4189 = new_n5534;
  assign po4190 = new_n5544;
  assign po4191 = new_n5545;
  assign po4192 = new_n5546;
  assign po4193 = new_n5547;
  assign po4194 = new_n5548;
  assign po4195 = new_n5549;
  assign po4196 = new_n5550;
  assign po4197 = new_n5551;
  assign po4198 = new_n5554;
  assign po4199 = new_n5555;
  assign po4200 = new_n5556;
  assign po4201 = new_n5557;
  assign po4202 = new_n5558;
  assign po4203 = new_n5559;
  assign po4204 = new_n5560;
  assign po4205 = new_n5561;
  assign po4206 = new_n5566;
  assign po4207 = new_n5567;
  assign po4208 = new_n5568;
  assign po4209 = new_n5569;
  assign po4210 = new_n5570;
  assign po4211 = new_n5571;
  assign po4212 = new_n5572;
  assign po4213 = new_n5573;
  assign po4214 = new_n5576;
  assign po4215 = new_n5577;
  assign po4216 = new_n5578;
  assign po4217 = new_n5579;
  assign po4218 = new_n5580;
  assign po4219 = new_n5581;
  assign po4220 = new_n5582;
  assign po4221 = new_n5583;
  assign po4222 = new_n5590;
  assign po4223 = new_n5591;
  assign po4224 = new_n5592;
  assign po4225 = new_n5593;
  assign po4226 = new_n5594;
  assign po4227 = new_n5595;
  assign po4228 = new_n5596;
  assign po4229 = new_n5597;
  assign po4230 = new_n5600;
  assign po4231 = new_n5601;
  assign po4232 = new_n5602;
  assign po4233 = new_n5603;
  assign po4234 = new_n5604;
  assign po4235 = new_n5605;
  assign po4236 = new_n5606;
  assign po4237 = new_n5607;
  assign po4238 = new_n5612;
  assign po4239 = new_n5613;
  assign po4240 = new_n5614;
  assign po4241 = new_n5615;
  assign po4242 = new_n5616;
  assign po4243 = new_n5617;
  assign po4244 = new_n5618;
  assign po4245 = new_n5619;
  assign po4246 = new_n5622;
  assign po4247 = new_n5623;
  assign po4248 = new_n5624;
  assign po4249 = new_n5625;
  assign po4250 = new_n5626;
  assign po4251 = new_n5627;
  assign po4252 = new_n5628;
  assign po4253 = new_n5629;
  assign po4254 = new_n5636;
  assign po4255 = new_n5637;
  assign po4256 = new_n5638;
  assign po4257 = new_n5639;
  assign po4258 = new_n5640;
  assign po4259 = new_n5641;
  assign po4260 = new_n5642;
  assign po4261 = new_n5643;
  assign po4262 = new_n5646;
  assign po4263 = new_n5647;
  assign po4264 = new_n5648;
  assign po4265 = new_n5649;
  assign po4266 = new_n5650;
  assign po4267 = new_n5651;
  assign po4268 = new_n5652;
  assign po4269 = new_n5653;
  assign po4270 = new_n5658;
  assign po4271 = new_n5659;
  assign po4272 = new_n5660;
  assign po4273 = new_n5661;
  assign po4274 = new_n5662;
  assign po4275 = new_n5663;
  assign po4276 = new_n5664;
  assign po4277 = new_n5665;
  assign po4278 = new_n5668;
  assign po4279 = new_n5669;
  assign po4280 = new_n5670;
  assign po4281 = new_n5671;
  assign po4282 = new_n5672;
  assign po4283 = new_n5673;
  assign po4284 = new_n5674;
  assign po4285 = new_n5675;
  assign po4286 = new_n5682;
  assign po4287 = new_n5683;
  assign po4288 = new_n5684;
  assign po4289 = new_n5685;
  assign po4290 = new_n5686;
  assign po4291 = new_n5687;
  assign po4292 = new_n5688;
  assign po4293 = new_n5689;
  assign po4294 = new_n5692;
  assign po4295 = new_n5693;
  assign po4296 = new_n5694;
  assign po4297 = new_n5695;
  assign po4298 = new_n5696;
  assign po4299 = new_n5697;
  assign po4300 = new_n5698;
  assign po4301 = new_n5699;
  assign po4302 = new_n5704;
  assign po4303 = new_n5705;
  assign po4304 = new_n5706;
  assign po4305 = new_n5707;
  assign po4306 = new_n5708;
  assign po4307 = new_n5709;
  assign po4308 = new_n5710;
  assign po4309 = new_n5711;
  assign po4310 = new_n5714;
  assign po4311 = new_n5715;
  assign po4312 = new_n5716;
  assign po4313 = new_n5717;
  assign po4314 = new_n5718;
  assign po4315 = new_n5719;
  assign po4316 = new_n5720;
  assign po4317 = new_n5721;
  assign po4318 = new_n5728;
  assign po4319 = new_n5729;
  assign po4320 = new_n5730;
  assign po4321 = new_n5731;
  assign po4322 = new_n5732;
  assign po4323 = new_n5733;
  assign po4324 = new_n5734;
  assign po4325 = new_n5735;
  assign po4326 = new_n5738;
  assign po4327 = new_n5739;
  assign po4328 = new_n5740;
  assign po4329 = new_n5741;
  assign po4330 = new_n5742;
  assign po4331 = new_n5743;
  assign po4332 = new_n5744;
  assign po4333 = new_n5745;
  assign po4334 = new_n5750;
  assign po4335 = new_n5751;
  assign po4336 = new_n5752;
  assign po4337 = new_n5753;
  assign po4338 = new_n5754;
  assign po4339 = new_n5755;
  assign po4340 = new_n5756;
  assign po4341 = new_n5757;
  assign po4342 = new_n5760;
  assign po4343 = new_n5761;
  assign po4344 = new_n5762;
  assign po4345 = new_n5763;
  assign po4346 = new_n5764;
  assign po4347 = new_n5765;
  assign po4348 = new_n5766;
  assign po4349 = new_n5767;
  assign po4350 = new_n5774;
  assign po4351 = new_n5775;
  assign po4352 = new_n5776;
  assign po4353 = new_n5777;
  assign po4354 = new_n5778;
  assign po4355 = new_n5779;
  assign po4356 = new_n5780;
  assign po4357 = new_n5781;
  assign po4358 = new_n5784;
  assign po4359 = new_n5785;
  assign po4360 = new_n5786;
  assign po4361 = new_n5787;
  assign po4362 = new_n5788;
  assign po4363 = new_n5789;
  assign po4364 = new_n5790;
  assign po4365 = new_n5791;
  assign po4366 = new_n5796;
  assign po4367 = new_n5797;
  assign po4368 = new_n5798;
  assign po4369 = new_n5799;
  assign po4370 = new_n5800;
  assign po4371 = new_n5801;
  assign po4372 = new_n5802;
  assign po4373 = new_n5803;
  assign po4374 = new_n5806;
  assign po4375 = new_n5807;
  assign po4376 = new_n5808;
  assign po4377 = new_n5809;
  assign po4378 = new_n5810;
  assign po4379 = new_n5811;
  assign po4380 = new_n5812;
  assign po4381 = new_n5813;
  assign po4382 = new_n5823;
  assign po4383 = new_n5824;
  assign po4384 = new_n5825;
  assign po4385 = new_n5826;
  assign po4386 = new_n5827;
  assign po4387 = new_n5828;
  assign po4388 = new_n5829;
  assign po4389 = new_n5830;
  assign po4390 = new_n5833;
  assign po4391 = new_n5834;
  assign po4392 = new_n5835;
  assign po4393 = new_n5836;
  assign po4394 = new_n5837;
  assign po4395 = new_n5838;
  assign po4396 = new_n5839;
  assign po4397 = new_n5840;
  assign po4398 = new_n5845;
  assign po4399 = new_n5846;
  assign po4400 = new_n5847;
  assign po4401 = new_n5848;
  assign po4402 = new_n5849;
  assign po4403 = new_n5850;
  assign po4404 = new_n5851;
  assign po4405 = new_n5852;
  assign po4406 = new_n5855;
  assign po4407 = new_n5856;
  assign po4408 = new_n5857;
  assign po4409 = new_n5858;
  assign po4410 = new_n5859;
  assign po4411 = new_n5860;
  assign po4412 = new_n5861;
  assign po4413 = new_n5862;
  assign po4414 = new_n5869;
  assign po4415 = new_n5870;
  assign po4416 = new_n5871;
  assign po4417 = new_n5872;
  assign po4418 = new_n5873;
  assign po4419 = new_n5874;
  assign po4420 = new_n5875;
  assign po4421 = new_n5876;
  assign po4422 = new_n5879;
  assign po4423 = new_n5880;
  assign po4424 = new_n5881;
  assign po4425 = new_n5882;
  assign po4426 = new_n5883;
  assign po4427 = new_n5884;
  assign po4428 = new_n5885;
  assign po4429 = new_n5886;
  assign po4430 = new_n5891;
  assign po4431 = new_n5892;
  assign po4432 = new_n5893;
  assign po4433 = new_n5894;
  assign po4434 = new_n5895;
  assign po4435 = new_n5896;
  assign po4436 = new_n5897;
  assign po4437 = new_n5898;
  assign po4438 = new_n5901;
  assign po4439 = new_n5902;
  assign po4440 = new_n5903;
  assign po4441 = new_n5904;
  assign po4442 = new_n5905;
  assign po4443 = new_n5906;
  assign po4444 = new_n5907;
  assign po4445 = new_n5908;
  assign po4446 = new_n5915;
  assign po4447 = new_n5916;
  assign po4448 = new_n5917;
  assign po4449 = new_n5918;
  assign po4450 = new_n5919;
  assign po4451 = new_n5920;
  assign po4452 = new_n5921;
  assign po4453 = new_n5922;
  assign po4454 = new_n5925;
  assign po4455 = new_n5926;
  assign po4456 = new_n5927;
  assign po4457 = new_n5928;
  assign po4458 = new_n5929;
  assign po4459 = new_n5930;
  assign po4460 = new_n5931;
  assign po4461 = new_n5932;
  assign po4462 = new_n5937;
  assign po4463 = new_n5938;
  assign po4464 = new_n5939;
  assign po4465 = new_n5940;
  assign po4466 = new_n5941;
  assign po4467 = new_n5942;
  assign po4468 = new_n5943;
  assign po4469 = new_n5944;
  assign po4470 = new_n5947;
  assign po4471 = new_n5948;
  assign po4472 = new_n5949;
  assign po4473 = new_n5950;
  assign po4474 = new_n5951;
  assign po4475 = new_n5952;
  assign po4476 = new_n5953;
  assign po4477 = new_n5954;
  assign po4478 = new_n5961;
  assign po4479 = new_n5962;
  assign po4480 = new_n5963;
  assign po4481 = new_n5964;
  assign po4482 = new_n5965;
  assign po4483 = new_n5966;
  assign po4484 = new_n5967;
  assign po4485 = new_n5968;
  assign po4486 = new_n5971;
  assign po4487 = new_n5972;
  assign po4488 = new_n5973;
  assign po4489 = new_n5974;
  assign po4490 = new_n5975;
  assign po4491 = new_n5976;
  assign po4492 = new_n5977;
  assign po4493 = new_n5978;
  assign po4494 = new_n5983;
  assign po4495 = new_n5984;
  assign po4496 = new_n5985;
  assign po4497 = new_n5986;
  assign po4498 = new_n5987;
  assign po4499 = new_n5988;
  assign po4500 = new_n5989;
  assign po4501 = new_n5990;
  assign po4502 = new_n5993;
  assign po4503 = new_n5994;
  assign po4504 = new_n5995;
  assign po4505 = new_n5996;
  assign po4506 = new_n5997;
  assign po4507 = new_n5998;
  assign po4508 = new_n5999;
  assign po4509 = new_n6000;
  assign po4510 = new_n6007;
  assign po4511 = new_n6008;
  assign po4512 = new_n6009;
  assign po4513 = new_n6010;
  assign po4514 = new_n6011;
  assign po4515 = new_n6012;
  assign po4516 = new_n6013;
  assign po4517 = new_n6014;
  assign po4518 = new_n6017;
  assign po4519 = new_n6018;
  assign po4520 = new_n6019;
  assign po4521 = new_n6020;
  assign po4522 = new_n6021;
  assign po4523 = new_n6022;
  assign po4524 = new_n6023;
  assign po4525 = new_n6024;
  assign po4526 = new_n6029;
  assign po4527 = new_n6030;
  assign po4528 = new_n6031;
  assign po4529 = new_n6032;
  assign po4530 = new_n6033;
  assign po4531 = new_n6034;
  assign po4532 = new_n6035;
  assign po4533 = new_n6036;
  assign po4534 = new_n6039;
  assign po4535 = new_n6040;
  assign po4536 = new_n6041;
  assign po4537 = new_n6042;
  assign po4538 = new_n6043;
  assign po4539 = new_n6044;
  assign po4540 = new_n6045;
  assign po4541 = new_n6046;
  assign po4542 = new_n6053;
  assign po4543 = new_n6054;
  assign po4544 = new_n6055;
  assign po4545 = new_n6056;
  assign po4546 = new_n6057;
  assign po4547 = new_n6058;
  assign po4548 = new_n6059;
  assign po4549 = new_n6060;
  assign po4550 = new_n6063;
  assign po4551 = new_n6064;
  assign po4552 = new_n6065;
  assign po4553 = new_n6066;
  assign po4554 = new_n6067;
  assign po4555 = new_n6068;
  assign po4556 = new_n6069;
  assign po4557 = new_n6070;
  assign po4558 = new_n6075;
  assign po4559 = new_n6076;
  assign po4560 = new_n6077;
  assign po4561 = new_n6078;
  assign po4562 = new_n6079;
  assign po4563 = new_n6080;
  assign po4564 = new_n6081;
  assign po4565 = new_n6082;
  assign po4566 = new_n6085;
  assign po4567 = new_n6086;
  assign po4568 = new_n6087;
  assign po4569 = new_n6088;
  assign po4570 = new_n6089;
  assign po4571 = new_n6090;
  assign po4572 = new_n6091;
  assign po4573 = new_n6092;
  assign po4574 = new_n6099;
  assign po4575 = new_n6100;
  assign po4576 = new_n6101;
  assign po4577 = new_n6102;
  assign po4578 = new_n6103;
  assign po4579 = new_n6104;
  assign po4580 = new_n6105;
  assign po4581 = new_n6106;
  assign po4582 = new_n6109;
  assign po4583 = new_n6110;
  assign po4584 = new_n6111;
  assign po4585 = new_n6112;
  assign po4586 = new_n6113;
  assign po4587 = new_n6114;
  assign po4588 = new_n6115;
  assign po4589 = new_n6116;
  assign po4590 = new_n6121;
  assign po4591 = new_n6122;
  assign po4592 = new_n6123;
  assign po4593 = new_n6124;
  assign po4594 = new_n6125;
  assign po4595 = new_n6126;
  assign po4596 = new_n6127;
  assign po4597 = new_n6128;
  assign po4598 = new_n6131;
  assign po4599 = new_n6132;
  assign po4600 = new_n6133;
  assign po4601 = new_n6134;
  assign po4602 = new_n6135;
  assign po4603 = new_n6136;
  assign po4604 = new_n6137;
  assign po4605 = new_n6138;
  assign po4606 = new_n6145;
  assign po4607 = new_n6146;
  assign po4608 = new_n6147;
  assign po4609 = new_n6148;
  assign po4610 = new_n6149;
  assign po4611 = new_n6150;
  assign po4612 = new_n6151;
  assign po4613 = new_n6152;
  assign po4614 = new_n6155;
  assign po4615 = new_n6156;
  assign po4616 = new_n6157;
  assign po4617 = new_n6158;
  assign po4618 = new_n6159;
  assign po4619 = new_n6160;
  assign po4620 = new_n6161;
  assign po4621 = new_n6162;
  assign po4622 = new_n6167;
  assign po4623 = new_n6168;
  assign po4624 = new_n6169;
  assign po4625 = new_n6170;
  assign po4626 = new_n6171;
  assign po4627 = new_n6172;
  assign po4628 = new_n6173;
  assign po4629 = new_n6174;
  assign po4630 = new_n6177;
  assign po4631 = new_n6178;
  assign po4632 = new_n6179;
  assign po4633 = new_n6180;
  assign po4634 = new_n6181;
  assign po4635 = new_n6182;
  assign po4636 = new_n6183;
  assign po4637 = new_n6184;
  assign po4638 = new_n6194;
  assign po4639 = new_n6195;
  assign po4640 = new_n6196;
  assign po4641 = new_n6197;
  assign po4642 = new_n6198;
  assign po4643 = new_n6199;
  assign po4644 = new_n6200;
  assign po4645 = new_n6201;
  assign po4646 = new_n6204;
  assign po4647 = new_n6205;
  assign po4648 = new_n6206;
  assign po4649 = new_n6207;
  assign po4650 = new_n6208;
  assign po4651 = new_n6209;
  assign po4652 = new_n6210;
  assign po4653 = new_n6211;
  assign po4654 = new_n6216;
  assign po4655 = new_n6217;
  assign po4656 = new_n6218;
  assign po4657 = new_n6219;
  assign po4658 = new_n6220;
  assign po4659 = new_n6221;
  assign po4660 = new_n6222;
  assign po4661 = new_n6223;
  assign po4662 = new_n6226;
  assign po4663 = new_n6227;
  assign po4664 = new_n6228;
  assign po4665 = new_n6229;
  assign po4666 = new_n6230;
  assign po4667 = new_n6231;
  assign po4668 = new_n6232;
  assign po4669 = new_n6233;
  assign po4670 = new_n6240;
  assign po4671 = new_n6241;
  assign po4672 = new_n6242;
  assign po4673 = new_n6243;
  assign po4674 = new_n6244;
  assign po4675 = new_n6245;
  assign po4676 = new_n6246;
  assign po4677 = new_n6247;
  assign po4678 = new_n6250;
  assign po4679 = new_n6251;
  assign po4680 = new_n6252;
  assign po4681 = new_n6253;
  assign po4682 = new_n6254;
  assign po4683 = new_n6255;
  assign po4684 = new_n6256;
  assign po4685 = new_n6257;
  assign po4686 = new_n6262;
  assign po4687 = new_n6263;
  assign po4688 = new_n6264;
  assign po4689 = new_n6265;
  assign po4690 = new_n6266;
  assign po4691 = new_n6267;
  assign po4692 = new_n6268;
  assign po4693 = new_n6269;
  assign po4694 = new_n6272;
  assign po4695 = new_n6273;
  assign po4696 = new_n6274;
  assign po4697 = new_n6275;
  assign po4698 = new_n6276;
  assign po4699 = new_n6277;
  assign po4700 = new_n6278;
  assign po4701 = new_n6279;
  assign po4702 = new_n6286;
  assign po4703 = new_n6287;
  assign po4704 = new_n6288;
  assign po4705 = new_n6289;
  assign po4706 = new_n6290;
  assign po4707 = new_n6291;
  assign po4708 = new_n6292;
  assign po4709 = new_n6293;
  assign po4710 = new_n6296;
  assign po4711 = new_n6297;
  assign po4712 = new_n6298;
  assign po4713 = new_n6299;
  assign po4714 = new_n6300;
  assign po4715 = new_n6301;
  assign po4716 = new_n6302;
  assign po4717 = new_n6303;
  assign po4718 = new_n6308;
  assign po4719 = new_n6309;
  assign po4720 = new_n6310;
  assign po4721 = new_n6311;
  assign po4722 = new_n6312;
  assign po4723 = new_n6313;
  assign po4724 = new_n6314;
  assign po4725 = new_n6315;
  assign po4726 = new_n6318;
  assign po4727 = new_n6319;
  assign po4728 = new_n6320;
  assign po4729 = new_n6321;
  assign po4730 = new_n6322;
  assign po4731 = new_n6323;
  assign po4732 = new_n6324;
  assign po4733 = new_n6325;
  assign po4734 = new_n6332;
  assign po4735 = new_n6333;
  assign po4736 = new_n6334;
  assign po4737 = new_n6335;
  assign po4738 = new_n6336;
  assign po4739 = new_n6337;
  assign po4740 = new_n6338;
  assign po4741 = new_n6339;
  assign po4742 = new_n6342;
  assign po4743 = new_n6343;
  assign po4744 = new_n6344;
  assign po4745 = new_n6345;
  assign po4746 = new_n6346;
  assign po4747 = new_n6347;
  assign po4748 = new_n6348;
  assign po4749 = new_n6349;
  assign po4750 = new_n6354;
  assign po4751 = new_n6355;
  assign po4752 = new_n6356;
  assign po4753 = new_n6357;
  assign po4754 = new_n6358;
  assign po4755 = new_n6359;
  assign po4756 = new_n6360;
  assign po4757 = new_n6361;
  assign po4758 = new_n6364;
  assign po4759 = new_n6365;
  assign po4760 = new_n6366;
  assign po4761 = new_n6367;
  assign po4762 = new_n6368;
  assign po4763 = new_n6369;
  assign po4764 = new_n6370;
  assign po4765 = new_n6371;
  assign po4766 = new_n6378;
  assign po4767 = new_n6379;
  assign po4768 = new_n6380;
  assign po4769 = new_n6381;
  assign po4770 = new_n6382;
  assign po4771 = new_n6383;
  assign po4772 = new_n6384;
  assign po4773 = new_n6385;
  assign po4774 = new_n6388;
  assign po4775 = new_n6389;
  assign po4776 = new_n6390;
  assign po4777 = new_n6391;
  assign po4778 = new_n6392;
  assign po4779 = new_n6393;
  assign po4780 = new_n6394;
  assign po4781 = new_n6395;
  assign po4782 = new_n6400;
  assign po4783 = new_n6401;
  assign po4784 = new_n6402;
  assign po4785 = new_n6403;
  assign po4786 = new_n6404;
  assign po4787 = new_n6405;
  assign po4788 = new_n6406;
  assign po4789 = new_n6407;
  assign po4790 = new_n6410;
  assign po4791 = new_n6411;
  assign po4792 = new_n6412;
  assign po4793 = new_n6413;
  assign po4794 = new_n6414;
  assign po4795 = new_n6415;
  assign po4796 = new_n6416;
  assign po4797 = new_n6417;
  assign po4798 = new_n6424;
  assign po4799 = new_n6425;
  assign po4800 = new_n6426;
  assign po4801 = new_n6427;
  assign po4802 = new_n6428;
  assign po4803 = new_n6429;
  assign po4804 = new_n6430;
  assign po4805 = new_n6431;
  assign po4806 = new_n6434;
  assign po4807 = new_n6435;
  assign po4808 = new_n6436;
  assign po4809 = new_n6437;
  assign po4810 = new_n6438;
  assign po4811 = new_n6439;
  assign po4812 = new_n6440;
  assign po4813 = new_n6441;
  assign po4814 = new_n6446;
  assign po4815 = new_n6447;
  assign po4816 = new_n6448;
  assign po4817 = new_n6449;
  assign po4818 = new_n6450;
  assign po4819 = new_n6451;
  assign po4820 = new_n6452;
  assign po4821 = new_n6453;
  assign po4822 = new_n6456;
  assign po4823 = new_n6457;
  assign po4824 = new_n6458;
  assign po4825 = new_n6459;
  assign po4826 = new_n6460;
  assign po4827 = new_n6461;
  assign po4828 = new_n6462;
  assign po4829 = new_n6463;
  assign po4830 = new_n6470;
  assign po4831 = new_n6471;
  assign po4832 = new_n6472;
  assign po4833 = new_n6473;
  assign po4834 = new_n6474;
  assign po4835 = new_n6475;
  assign po4836 = new_n6476;
  assign po4837 = new_n6477;
  assign po4838 = new_n6480;
  assign po4839 = new_n6481;
  assign po4840 = new_n6482;
  assign po4841 = new_n6483;
  assign po4842 = new_n6484;
  assign po4843 = new_n6485;
  assign po4844 = new_n6486;
  assign po4845 = new_n6487;
  assign po4846 = new_n6492;
  assign po4847 = new_n6493;
  assign po4848 = new_n6494;
  assign po4849 = new_n6495;
  assign po4850 = new_n6496;
  assign po4851 = new_n6497;
  assign po4852 = new_n6498;
  assign po4853 = new_n6499;
  assign po4854 = new_n6502;
  assign po4855 = new_n6503;
  assign po4856 = new_n6504;
  assign po4857 = new_n6505;
  assign po4858 = new_n6506;
  assign po4859 = new_n6507;
  assign po4860 = new_n6508;
  assign po4861 = new_n6509;
  assign po4862 = new_n6516;
  assign po4863 = new_n6517;
  assign po4864 = new_n6518;
  assign po4865 = new_n6519;
  assign po4866 = new_n6520;
  assign po4867 = new_n6521;
  assign po4868 = new_n6522;
  assign po4869 = new_n6523;
  assign po4870 = new_n6526;
  assign po4871 = new_n6527;
  assign po4872 = new_n6528;
  assign po4873 = new_n6529;
  assign po4874 = new_n6530;
  assign po4875 = new_n6531;
  assign po4876 = new_n6532;
  assign po4877 = new_n6533;
  assign po4878 = new_n6538;
  assign po4879 = new_n6539;
  assign po4880 = new_n6540;
  assign po4881 = new_n6541;
  assign po4882 = new_n6542;
  assign po4883 = new_n6543;
  assign po4884 = new_n6544;
  assign po4885 = new_n6545;
  assign po4886 = new_n6548;
  assign po4887 = new_n6549;
  assign po4888 = new_n6550;
  assign po4889 = new_n6551;
  assign po4890 = new_n6552;
  assign po4891 = new_n6553;
  assign po4892 = new_n6554;
  assign po4893 = new_n6555;
  assign po4894 = new_n6565;
  assign po4895 = new_n6566;
  assign po4896 = new_n6567;
  assign po4897 = new_n6568;
  assign po4898 = new_n6569;
  assign po4899 = new_n6570;
  assign po4900 = new_n6571;
  assign po4901 = new_n6572;
  assign po4902 = new_n6575;
  assign po4903 = new_n6576;
  assign po4904 = new_n6577;
  assign po4905 = new_n6578;
  assign po4906 = new_n6579;
  assign po4907 = new_n6580;
  assign po4908 = new_n6581;
  assign po4909 = new_n6582;
  assign po4910 = new_n6587;
  assign po4911 = new_n6588;
  assign po4912 = new_n6589;
  assign po4913 = new_n6590;
  assign po4914 = new_n6591;
  assign po4915 = new_n6592;
  assign po4916 = new_n6593;
  assign po4917 = new_n6594;
  assign po4918 = new_n6597;
  assign po4919 = new_n6598;
  assign po4920 = new_n6599;
  assign po4921 = new_n6600;
  assign po4922 = new_n6601;
  assign po4923 = new_n6602;
  assign po4924 = new_n6603;
  assign po4925 = new_n6604;
  assign po4926 = new_n6611;
  assign po4927 = new_n6612;
  assign po4928 = new_n6613;
  assign po4929 = new_n6614;
  assign po4930 = new_n6615;
  assign po4931 = new_n6616;
  assign po4932 = new_n6617;
  assign po4933 = new_n6618;
  assign po4934 = new_n6621;
  assign po4935 = new_n6622;
  assign po4936 = new_n6623;
  assign po4937 = new_n6624;
  assign po4938 = new_n6625;
  assign po4939 = new_n6626;
  assign po4940 = new_n6627;
  assign po4941 = new_n6628;
  assign po4942 = new_n6633;
  assign po4943 = new_n6634;
  assign po4944 = new_n6635;
  assign po4945 = new_n6636;
  assign po4946 = new_n6637;
  assign po4947 = new_n6638;
  assign po4948 = new_n6639;
  assign po4949 = new_n6640;
  assign po4950 = new_n6643;
  assign po4951 = new_n6644;
  assign po4952 = new_n6645;
  assign po4953 = new_n6646;
  assign po4954 = new_n6647;
  assign po4955 = new_n6648;
  assign po4956 = new_n6649;
  assign po4957 = new_n6650;
  assign po4958 = new_n6657;
  assign po4959 = new_n6658;
  assign po4960 = new_n6659;
  assign po4961 = new_n6660;
  assign po4962 = new_n6661;
  assign po4963 = new_n6662;
  assign po4964 = new_n6663;
  assign po4965 = new_n6664;
  assign po4966 = new_n6667;
  assign po4967 = new_n6668;
  assign po4968 = new_n6669;
  assign po4969 = new_n6670;
  assign po4970 = new_n6671;
  assign po4971 = new_n6672;
  assign po4972 = new_n6673;
  assign po4973 = new_n6674;
  assign po4974 = new_n6679;
  assign po4975 = new_n6680;
  assign po4976 = new_n6681;
  assign po4977 = new_n6682;
  assign po4978 = new_n6683;
  assign po4979 = new_n6684;
  assign po4980 = new_n6685;
  assign po4981 = new_n6686;
  assign po4982 = new_n6689;
  assign po4983 = new_n6690;
  assign po4984 = new_n6691;
  assign po4985 = new_n6692;
  assign po4986 = new_n6693;
  assign po4987 = new_n6694;
  assign po4988 = new_n6695;
  assign po4989 = new_n6696;
  assign po4990 = new_n6703;
  assign po4991 = new_n6704;
  assign po4992 = new_n6705;
  assign po4993 = new_n6706;
  assign po4994 = new_n6707;
  assign po4995 = new_n6708;
  assign po4996 = new_n6709;
  assign po4997 = new_n6710;
  assign po4998 = new_n6713;
  assign po4999 = new_n6714;
  assign po5000 = new_n6715;
  assign po5001 = new_n6716;
  assign po5002 = new_n6717;
  assign po5003 = new_n6718;
  assign po5004 = new_n6719;
  assign po5005 = new_n6720;
  assign po5006 = new_n6725;
  assign po5007 = new_n6726;
  assign po5008 = new_n6727;
  assign po5009 = new_n6728;
  assign po5010 = new_n6729;
  assign po5011 = new_n6730;
  assign po5012 = new_n6731;
  assign po5013 = new_n6732;
  assign po5014 = new_n6735;
  assign po5015 = new_n6736;
  assign po5016 = new_n6737;
  assign po5017 = new_n6738;
  assign po5018 = new_n6739;
  assign po5019 = new_n6740;
  assign po5020 = new_n6741;
  assign po5021 = new_n6742;
  assign po5022 = new_n6749;
  assign po5023 = new_n6750;
  assign po5024 = new_n6751;
  assign po5025 = new_n6752;
  assign po5026 = new_n6753;
  assign po5027 = new_n6754;
  assign po5028 = new_n6755;
  assign po5029 = new_n6756;
  assign po5030 = new_n6759;
  assign po5031 = new_n6760;
  assign po5032 = new_n6761;
  assign po5033 = new_n6762;
  assign po5034 = new_n6763;
  assign po5035 = new_n6764;
  assign po5036 = new_n6765;
  assign po5037 = new_n6766;
  assign po5038 = new_n6771;
  assign po5039 = new_n6772;
  assign po5040 = new_n6773;
  assign po5041 = new_n6774;
  assign po5042 = new_n6775;
  assign po5043 = new_n6776;
  assign po5044 = new_n6777;
  assign po5045 = new_n6778;
  assign po5046 = new_n6781;
  assign po5047 = new_n6782;
  assign po5048 = new_n6783;
  assign po5049 = new_n6784;
  assign po5050 = new_n6785;
  assign po5051 = new_n6786;
  assign po5052 = new_n6787;
  assign po5053 = new_n6788;
  assign po5054 = new_n6795;
  assign po5055 = new_n6796;
  assign po5056 = new_n6797;
  assign po5057 = new_n6798;
  assign po5058 = new_n6799;
  assign po5059 = new_n6800;
  assign po5060 = new_n6801;
  assign po5061 = new_n6802;
  assign po5062 = new_n6805;
  assign po5063 = new_n6806;
  assign po5064 = new_n6807;
  assign po5065 = new_n6808;
  assign po5066 = new_n6809;
  assign po5067 = new_n6810;
  assign po5068 = new_n6811;
  assign po5069 = new_n6812;
  assign po5070 = new_n6817;
  assign po5071 = new_n6818;
  assign po5072 = new_n6819;
  assign po5073 = new_n6820;
  assign po5074 = new_n6821;
  assign po5075 = new_n6822;
  assign po5076 = new_n6823;
  assign po5077 = new_n6824;
  assign po5078 = new_n6827;
  assign po5079 = new_n6828;
  assign po5080 = new_n6829;
  assign po5081 = new_n6830;
  assign po5082 = new_n6831;
  assign po5083 = new_n6832;
  assign po5084 = new_n6833;
  assign po5085 = new_n6834;
  assign po5086 = new_n6841;
  assign po5087 = new_n6842;
  assign po5088 = new_n6843;
  assign po5089 = new_n6844;
  assign po5090 = new_n6845;
  assign po5091 = new_n6846;
  assign po5092 = new_n6847;
  assign po5093 = new_n6848;
  assign po5094 = new_n6851;
  assign po5095 = new_n6852;
  assign po5096 = new_n6853;
  assign po5097 = new_n6854;
  assign po5098 = new_n6855;
  assign po5099 = new_n6856;
  assign po5100 = new_n6857;
  assign po5101 = new_n6858;
  assign po5102 = new_n6863;
  assign po5103 = new_n6864;
  assign po5104 = new_n6865;
  assign po5105 = new_n6866;
  assign po5106 = new_n6867;
  assign po5107 = new_n6868;
  assign po5108 = new_n6869;
  assign po5109 = new_n6870;
  assign po5110 = new_n6873;
  assign po5111 = new_n6874;
  assign po5112 = new_n6875;
  assign po5113 = new_n6876;
  assign po5114 = new_n6877;
  assign po5115 = new_n6878;
  assign po5116 = new_n6879;
  assign po5117 = new_n6880;
  assign po5118 = new_n6887;
  assign po5119 = new_n6888;
  assign po5120 = new_n6889;
  assign po5121 = new_n6890;
  assign po5122 = new_n6891;
  assign po5123 = new_n6892;
  assign po5124 = new_n6893;
  assign po5125 = new_n6894;
  assign po5126 = new_n6897;
  assign po5127 = new_n6898;
  assign po5128 = new_n6899;
  assign po5129 = new_n6900;
  assign po5130 = new_n6901;
  assign po5131 = new_n6902;
  assign po5132 = new_n6903;
  assign po5133 = new_n6904;
  assign po5134 = new_n6909;
  assign po5135 = new_n6910;
  assign po5136 = new_n6911;
  assign po5137 = new_n6912;
  assign po5138 = new_n6913;
  assign po5139 = new_n6914;
  assign po5140 = new_n6915;
  assign po5141 = new_n6916;
  assign po5142 = new_n6919;
  assign po5143 = new_n6920;
  assign po5144 = new_n6921;
  assign po5145 = new_n6922;
  assign po5146 = new_n6923;
  assign po5147 = new_n6924;
  assign po5148 = new_n6925;
  assign po5149 = new_n6926;
  assign po5150 = new_n6933;
  assign po5151 = new_n6934;
  assign po5152 = new_n6935;
  assign po5153 = new_n6936;
  assign po5154 = new_n6937;
  assign po5155 = new_n6938;
  assign po5156 = new_n6939;
  assign po5157 = new_n6940;
  assign po5158 = new_n6943;
  assign po5159 = new_n6944;
  assign po5160 = new_n6945;
  assign po5161 = new_n6946;
  assign po5162 = new_n6947;
  assign po5163 = new_n6948;
  assign po5164 = new_n6949;
  assign po5165 = new_n6950;
  assign po5166 = new_n6955;
  assign po5167 = new_n6956;
  assign po5168 = new_n6957;
  assign po5169 = new_n6958;
  assign po5170 = new_n6959;
  assign po5171 = new_n6960;
  assign po5172 = new_n6961;
  assign po5173 = new_n6962;
  assign po5174 = new_n6965;
  assign po5175 = new_n6966;
  assign po5176 = new_n6967;
  assign po5177 = new_n6968;
  assign po5178 = new_n6969;
  assign po5179 = new_n6970;
  assign po5180 = new_n6971;
  assign po5181 = new_n6972;
  assign po5182 = new_n6979;
  assign po5183 = new_n6980;
  assign po5184 = new_n6981;
  assign po5185 = new_n6982;
  assign po5186 = new_n6983;
  assign po5187 = new_n6984;
  assign po5188 = new_n6985;
  assign po5189 = new_n6986;
  assign po5190 = new_n6989;
  assign po5191 = new_n6990;
  assign po5192 = new_n6991;
  assign po5193 = new_n6992;
  assign po5194 = new_n6993;
  assign po5195 = new_n6994;
  assign po5196 = new_n6995;
  assign po5197 = new_n6996;
  assign po5198 = new_n7001;
  assign po5199 = new_n7002;
  assign po5200 = new_n7003;
  assign po5201 = new_n7004;
  assign po5202 = new_n7005;
  assign po5203 = new_n7006;
  assign po5204 = new_n7007;
  assign po5205 = new_n7008;
  assign po5206 = new_n7011;
  assign po5207 = new_n7012;
  assign po5208 = new_n7013;
  assign po5209 = new_n7014;
  assign po5210 = new_n7015;
  assign po5211 = new_n7016;
  assign po5212 = new_n7017;
  assign po5213 = new_n7018;
  assign po5214 = new_n7025;
  assign po5215 = new_n7026;
  assign po5216 = new_n7027;
  assign po5217 = new_n7028;
  assign po5218 = new_n7029;
  assign po5219 = new_n7030;
  assign po5220 = new_n7031;
  assign po5221 = new_n7032;
  assign po5222 = new_n7035;
  assign po5223 = new_n7036;
  assign po5224 = new_n7037;
  assign po5225 = new_n7038;
  assign po5226 = new_n7039;
  assign po5227 = new_n7040;
  assign po5228 = new_n7041;
  assign po5229 = new_n7042;
  assign po5230 = new_n7047;
  assign po5231 = new_n7048;
  assign po5232 = new_n7049;
  assign po5233 = new_n7050;
  assign po5234 = new_n7051;
  assign po5235 = new_n7052;
  assign po5236 = new_n7053;
  assign po5237 = new_n7054;
  assign po5238 = new_n7057;
  assign po5239 = new_n7058;
  assign po5240 = new_n7059;
  assign po5241 = new_n7060;
  assign po5242 = new_n7061;
  assign po5243 = new_n7062;
  assign po5244 = new_n7063;
  assign po5245 = new_n7064;
  assign po5246 = new_n7071;
  assign po5247 = new_n7072;
  assign po5248 = new_n7073;
  assign po5249 = new_n7074;
  assign po5250 = new_n7075;
  assign po5251 = new_n7076;
  assign po5252 = new_n7077;
  assign po5253 = new_n7078;
  assign po5254 = new_n7081;
  assign po5255 = new_n7082;
  assign po5256 = new_n7083;
  assign po5257 = new_n7084;
  assign po5258 = new_n7085;
  assign po5259 = new_n7086;
  assign po5260 = new_n7087;
  assign po5261 = new_n7088;
  assign po5262 = new_n7093;
  assign po5263 = new_n7094;
  assign po5264 = new_n7095;
  assign po5265 = new_n7096;
  assign po5266 = new_n7097;
  assign po5267 = new_n7098;
  assign po5268 = new_n7099;
  assign po5269 = new_n7100;
  assign po5270 = new_n7103;
  assign po5271 = new_n7104;
  assign po5272 = new_n7105;
  assign po5273 = new_n7106;
  assign po5274 = new_n7107;
  assign po5275 = new_n7108;
  assign po5276 = new_n7109;
  assign po5277 = new_n7110;
  assign po5278 = new_n7117;
  assign po5279 = new_n7118;
  assign po5280 = new_n7119;
  assign po5281 = new_n7120;
  assign po5282 = new_n7121;
  assign po5283 = new_n7122;
  assign po5284 = new_n7123;
  assign po5285 = new_n7124;
  assign po5286 = new_n7127;
  assign po5287 = new_n7128;
  assign po5288 = new_n7129;
  assign po5289 = new_n7130;
  assign po5290 = new_n7131;
  assign po5291 = new_n7132;
  assign po5292 = new_n7133;
  assign po5293 = new_n7134;
  assign po5294 = new_n7139;
  assign po5295 = new_n7140;
  assign po5296 = new_n7141;
  assign po5297 = new_n7142;
  assign po5298 = new_n7143;
  assign po5299 = new_n7144;
  assign po5300 = new_n7145;
  assign po5301 = new_n7146;
  assign po5302 = new_n7149;
  assign po5303 = new_n7150;
  assign po5304 = new_n7151;
  assign po5305 = new_n7152;
  assign po5306 = new_n7153;
  assign po5307 = new_n7154;
  assign po5308 = new_n7155;
  assign po5309 = new_n7156;
  assign po5310 = new_n7163;
  assign po5311 = new_n7164;
  assign po5312 = new_n7165;
  assign po5313 = new_n7166;
  assign po5314 = new_n7167;
  assign po5315 = new_n7168;
  assign po5316 = new_n7169;
  assign po5317 = new_n7170;
  assign po5318 = new_n7173;
  assign po5319 = new_n7174;
  assign po5320 = new_n7175;
  assign po5321 = new_n7176;
  assign po5322 = new_n7177;
  assign po5323 = new_n7178;
  assign po5324 = new_n7179;
  assign po5325 = new_n7180;
  assign po5326 = new_n7185;
  assign po5327 = new_n7186;
  assign po5328 = new_n7187;
  assign po5329 = new_n7188;
  assign po5330 = new_n7189;
  assign po5331 = new_n7190;
  assign po5332 = new_n7191;
  assign po5333 = new_n7192;
  assign po5334 = new_n7195;
  assign po5335 = new_n7196;
  assign po5336 = new_n7197;
  assign po5337 = new_n7198;
  assign po5338 = new_n7199;
  assign po5339 = new_n7200;
  assign po5340 = new_n7201;
  assign po5341 = new_n7202;
  assign po5342 = new_n7209;
  assign po5343 = new_n7210;
  assign po5344 = new_n7211;
  assign po5345 = new_n7212;
  assign po5346 = new_n7213;
  assign po5347 = new_n7214;
  assign po5348 = new_n7215;
  assign po5349 = new_n7216;
  assign po5350 = new_n7219;
  assign po5351 = new_n7220;
  assign po5352 = new_n7221;
  assign po5353 = new_n7222;
  assign po5354 = new_n7223;
  assign po5355 = new_n7224;
  assign po5356 = new_n7225;
  assign po5357 = new_n7226;
  assign po5358 = new_n7231;
  assign po5359 = new_n7232;
  assign po5360 = new_n7233;
  assign po5361 = new_n7234;
  assign po5362 = new_n7235;
  assign po5363 = new_n7236;
  assign po5364 = new_n7237;
  assign po5365 = new_n7238;
  assign po5366 = new_n7241;
  assign po5367 = new_n7242;
  assign po5368 = new_n7243;
  assign po5369 = new_n7244;
  assign po5370 = new_n7245;
  assign po5371 = new_n7246;
  assign po5372 = new_n7247;
  assign po5373 = new_n7248;
  assign po5374 = new_n7255;
  assign po5375 = new_n7256;
  assign po5376 = new_n7257;
  assign po5377 = new_n7258;
  assign po5378 = new_n7259;
  assign po5379 = new_n7260;
  assign po5380 = new_n7261;
  assign po5381 = new_n7262;
  assign po5382 = new_n7265;
  assign po5383 = new_n7266;
  assign po5384 = new_n7267;
  assign po5385 = new_n7268;
  assign po5386 = new_n7269;
  assign po5387 = new_n7270;
  assign po5388 = new_n7271;
  assign po5389 = new_n7272;
  assign po5390 = new_n7277;
  assign po5391 = new_n7278;
  assign po5392 = new_n7279;
  assign po5393 = new_n7280;
  assign po5394 = new_n7281;
  assign po5395 = new_n7282;
  assign po5396 = new_n7283;
  assign po5397 = new_n7284;
  assign po5398 = new_n7287;
  assign po5399 = new_n7288;
  assign po5400 = new_n7289;
  assign po5401 = new_n7290;
  assign po5402 = new_n7291;
  assign po5403 = new_n7292;
  assign po5404 = new_n7293;
  assign po5405 = new_n7294;
  assign po5406 = new_n7301;
  assign po5407 = new_n7302;
  assign po5408 = new_n7303;
  assign po5409 = new_n7304;
  assign po5410 = new_n7305;
  assign po5411 = new_n7306;
  assign po5412 = new_n7307;
  assign po5413 = new_n7308;
  assign po5414 = new_n7311;
  assign po5415 = new_n7312;
  assign po5416 = new_n7313;
  assign po5417 = new_n7314;
  assign po5418 = new_n7315;
  assign po5419 = new_n7316;
  assign po5420 = new_n7317;
  assign po5421 = new_n7318;
  assign po5422 = new_n7323;
  assign po5423 = new_n7324;
  assign po5424 = new_n7325;
  assign po5425 = new_n7326;
  assign po5426 = new_n7327;
  assign po5427 = new_n7328;
  assign po5428 = new_n7329;
  assign po5429 = new_n7330;
  assign po5430 = new_n7333;
  assign po5431 = new_n7334;
  assign po5432 = new_n7335;
  assign po5433 = new_n7336;
  assign po5434 = new_n7337;
  assign po5435 = new_n7338;
  assign po5436 = new_n7339;
  assign po5437 = new_n7340;
  assign po5438 = new_n7347;
  assign po5439 = new_n7348;
  assign po5440 = new_n7349;
  assign po5441 = new_n7350;
  assign po5442 = new_n7351;
  assign po5443 = new_n7352;
  assign po5444 = new_n7353;
  assign po5445 = new_n7354;
  assign po5446 = new_n7357;
  assign po5447 = new_n7358;
  assign po5448 = new_n7359;
  assign po5449 = new_n7360;
  assign po5450 = new_n7361;
  assign po5451 = new_n7362;
  assign po5452 = new_n7363;
  assign po5453 = new_n7364;
  assign po5454 = new_n7369;
  assign po5455 = new_n7370;
  assign po5456 = new_n7371;
  assign po5457 = new_n7372;
  assign po5458 = new_n7373;
  assign po5459 = new_n7374;
  assign po5460 = new_n7375;
  assign po5461 = new_n7376;
  assign po5462 = new_n7379;
  assign po5463 = new_n7380;
  assign po5464 = new_n7381;
  assign po5465 = new_n7382;
  assign po5466 = new_n7383;
  assign po5467 = new_n7384;
  assign po5468 = new_n7385;
  assign po5469 = new_n7386;
  assign po5470 = new_n7393;
  assign po5471 = new_n7394;
  assign po5472 = new_n7395;
  assign po5473 = new_n7396;
  assign po5474 = new_n7397;
  assign po5475 = new_n7398;
  assign po5476 = new_n7399;
  assign po5477 = new_n7400;
  assign po5478 = new_n7403;
  assign po5479 = new_n7404;
  assign po5480 = new_n7405;
  assign po5481 = new_n7406;
  assign po5482 = new_n7407;
  assign po5483 = new_n7408;
  assign po5484 = new_n7409;
  assign po5485 = new_n7410;
  assign po5486 = new_n7415;
  assign po5487 = new_n7416;
  assign po5488 = new_n7417;
  assign po5489 = new_n7418;
  assign po5490 = new_n7419;
  assign po5491 = new_n7420;
  assign po5492 = new_n7421;
  assign po5493 = new_n7422;
  assign po5494 = new_n7425;
  assign po5495 = new_n7426;
  assign po5496 = new_n7427;
  assign po5497 = new_n7428;
  assign po5498 = new_n7429;
  assign po5499 = new_n7430;
  assign po5500 = new_n7431;
  assign po5501 = new_n7432;
  assign po5502 = new_n7439;
  assign po5503 = new_n7440;
  assign po5504 = new_n7441;
  assign po5505 = new_n7442;
  assign po5506 = new_n7443;
  assign po5507 = new_n7444;
  assign po5508 = new_n7445;
  assign po5509 = new_n7446;
  assign po5510 = new_n7449;
  assign po5511 = new_n7450;
  assign po5512 = new_n7451;
  assign po5513 = new_n7452;
  assign po5514 = new_n7453;
  assign po5515 = new_n7454;
  assign po5516 = new_n7455;
  assign po5517 = new_n7456;
  assign po5518 = new_n7461;
  assign po5519 = new_n7462;
  assign po5520 = new_n7463;
  assign po5521 = new_n7464;
  assign po5522 = new_n7465;
  assign po5523 = new_n7466;
  assign po5524 = new_n7467;
  assign po5525 = new_n7468;
  assign po5526 = new_n7471;
  assign po5527 = new_n7472;
  assign po5528 = new_n7473;
  assign po5529 = new_n7474;
  assign po5530 = new_n7475;
  assign po5531 = new_n7476;
  assign po5532 = new_n7477;
  assign po5533 = new_n7478;
  assign po5534 = new_n7485;
  assign po5535 = new_n7486;
  assign po5536 = new_n7487;
  assign po5537 = new_n7488;
  assign po5538 = new_n7489;
  assign po5539 = new_n7490;
  assign po5540 = new_n7491;
  assign po5541 = new_n7492;
  assign po5542 = new_n7495;
  assign po5543 = new_n7496;
  assign po5544 = new_n7497;
  assign po5545 = new_n7498;
  assign po5546 = new_n7499;
  assign po5547 = new_n7500;
  assign po5548 = new_n7501;
  assign po5549 = new_n7502;
  assign po5550 = new_n7507;
  assign po5551 = new_n7508;
  assign po5552 = new_n7509;
  assign po5553 = new_n7510;
  assign po5554 = new_n7511;
  assign po5555 = new_n7512;
  assign po5556 = new_n7513;
  assign po5557 = new_n7514;
  assign po5558 = new_n7517;
  assign po5559 = new_n7518;
  assign po5560 = new_n7519;
  assign po5561 = new_n7520;
  assign po5562 = new_n7521;
  assign po5563 = new_n7522;
  assign po5564 = new_n7523;
  assign po5565 = new_n7524;
  assign po5566 = new_n7531;
  assign po5567 = new_n7532;
  assign po5568 = new_n7533;
  assign po5569 = new_n7534;
  assign po5570 = new_n7535;
  assign po5571 = new_n7536;
  assign po5572 = new_n7537;
  assign po5573 = new_n7538;
  assign po5574 = new_n7541;
  assign po5575 = new_n7542;
  assign po5576 = new_n7543;
  assign po5577 = new_n7544;
  assign po5578 = new_n7545;
  assign po5579 = new_n7546;
  assign po5580 = new_n7547;
  assign po5581 = new_n7548;
  assign po5582 = new_n7553;
  assign po5583 = new_n7554;
  assign po5584 = new_n7555;
  assign po5585 = new_n7556;
  assign po5586 = new_n7557;
  assign po5587 = new_n7558;
  assign po5588 = new_n7559;
  assign po5589 = new_n7560;
  assign po5590 = new_n7563;
  assign po5591 = new_n7564;
  assign po5592 = new_n7565;
  assign po5593 = new_n7566;
  assign po5594 = new_n7567;
  assign po5595 = new_n7568;
  assign po5596 = new_n7569;
  assign po5597 = new_n7570;
  assign po5598 = new_n7577;
  assign po5599 = new_n7578;
  assign po5600 = new_n7579;
  assign po5601 = new_n7580;
  assign po5602 = new_n7581;
  assign po5603 = new_n7582;
  assign po5604 = new_n7583;
  assign po5605 = new_n7584;
  assign po5606 = new_n7587;
  assign po5607 = new_n7588;
  assign po5608 = new_n7589;
  assign po5609 = new_n7590;
  assign po5610 = new_n7591;
  assign po5611 = new_n7592;
  assign po5612 = new_n7593;
  assign po5613 = new_n7594;
  assign po5614 = new_n7599;
  assign po5615 = new_n7600;
  assign po5616 = new_n7601;
  assign po5617 = new_n7602;
  assign po5618 = new_n7603;
  assign po5619 = new_n7604;
  assign po5620 = new_n7605;
  assign po5621 = new_n7606;
  assign po5622 = new_n7609;
  assign po5623 = new_n7610;
  assign po5624 = new_n7611;
  assign po5625 = new_n7612;
  assign po5626 = new_n7613;
  assign po5627 = new_n7614;
  assign po5628 = new_n7615;
  assign po5629 = new_n7616;
  assign po5630 = new_n7623;
  assign po5631 = new_n7624;
  assign po5632 = new_n7625;
  assign po5633 = new_n7626;
  assign po5634 = new_n7627;
  assign po5635 = new_n7628;
  assign po5636 = new_n7629;
  assign po5637 = new_n7630;
  assign po5638 = new_n7633;
  assign po5639 = new_n7634;
  assign po5640 = new_n7635;
  assign po5641 = new_n7636;
  assign po5642 = new_n7637;
  assign po5643 = new_n7638;
  assign po5644 = new_n7639;
  assign po5645 = new_n7640;
  assign po5646 = new_n7645;
  assign po5647 = new_n7646;
  assign po5648 = new_n7647;
  assign po5649 = new_n7648;
  assign po5650 = new_n7649;
  assign po5651 = new_n7650;
  assign po5652 = new_n7651;
  assign po5653 = new_n7652;
  assign po5654 = new_n7655;
  assign po5655 = new_n7656;
  assign po5656 = new_n7657;
  assign po5657 = new_n7658;
  assign po5658 = new_n7659;
  assign po5659 = new_n7660;
  assign po5660 = new_n7661;
  assign po5661 = new_n7662;
  assign po5662 = new_n7669;
  assign po5663 = new_n7670;
  assign po5664 = new_n7671;
  assign po5665 = new_n7672;
  assign po5666 = new_n7673;
  assign po5667 = new_n7674;
  assign po5668 = new_n7675;
  assign po5669 = new_n7676;
  assign po5670 = new_n7679;
  assign po5671 = new_n7680;
  assign po5672 = new_n7681;
  assign po5673 = new_n7682;
  assign po5674 = new_n7683;
  assign po5675 = new_n7684;
  assign po5676 = new_n7685;
  assign po5677 = new_n7686;
  assign po5678 = new_n7691;
  assign po5679 = new_n7692;
  assign po5680 = new_n7693;
  assign po5681 = new_n7694;
  assign po5682 = new_n7695;
  assign po5683 = new_n7696;
  assign po5684 = new_n7697;
  assign po5685 = new_n7698;
  assign po5686 = new_n7701;
  assign po5687 = new_n7702;
  assign po5688 = new_n7703;
  assign po5689 = new_n7704;
  assign po5690 = new_n7705;
  assign po5691 = new_n7706;
  assign po5692 = new_n7707;
  assign po5693 = new_n7708;
  assign po5694 = new_n7715;
  assign po5695 = new_n7716;
  assign po5696 = new_n7717;
  assign po5697 = new_n7718;
  assign po5698 = new_n7719;
  assign po5699 = new_n7720;
  assign po5700 = new_n7721;
  assign po5701 = new_n7722;
  assign po5702 = new_n7725;
  assign po5703 = new_n7726;
  assign po5704 = new_n7727;
  assign po5705 = new_n7728;
  assign po5706 = new_n7729;
  assign po5707 = new_n7730;
  assign po5708 = new_n7731;
  assign po5709 = new_n7732;
  assign po5710 = new_n7737;
  assign po5711 = new_n7738;
  assign po5712 = new_n7739;
  assign po5713 = new_n7740;
  assign po5714 = new_n7741;
  assign po5715 = new_n7742;
  assign po5716 = new_n7743;
  assign po5717 = new_n7744;
  assign po5718 = new_n7747;
  assign po5719 = new_n7748;
  assign po5720 = new_n7749;
  assign po5721 = new_n7750;
  assign po5722 = new_n7751;
  assign po5723 = new_n7752;
  assign po5724 = new_n7753;
  assign po5725 = new_n7754;
  assign po5726 = new_n7761;
  assign po5727 = new_n7762;
  assign po5728 = new_n7763;
  assign po5729 = new_n7764;
  assign po5730 = new_n7765;
  assign po5731 = new_n7766;
  assign po5732 = new_n7767;
  assign po5733 = new_n7768;
  assign po5734 = new_n7771;
  assign po5735 = new_n7772;
  assign po5736 = new_n7773;
  assign po5737 = new_n7774;
  assign po5738 = new_n7775;
  assign po5739 = new_n7776;
  assign po5740 = new_n7777;
  assign po5741 = new_n7778;
  assign po5742 = new_n7783;
  assign po5743 = new_n7784;
  assign po5744 = new_n7785;
  assign po5745 = new_n7786;
  assign po5746 = new_n7787;
  assign po5747 = new_n7788;
  assign po5748 = new_n7789;
  assign po5749 = new_n7790;
  assign po5750 = new_n7793;
  assign po5751 = new_n7794;
  assign po5752 = new_n7795;
  assign po5753 = new_n7796;
  assign po5754 = new_n7797;
  assign po5755 = new_n7798;
  assign po5756 = new_n7799;
  assign po5757 = new_n7800;
  assign po5758 = new_n7807;
  assign po5759 = new_n7808;
  assign po5760 = new_n7809;
  assign po5761 = new_n7810;
  assign po5762 = new_n7811;
  assign po5763 = new_n7812;
  assign po5764 = new_n7813;
  assign po5765 = new_n7814;
  assign po5766 = new_n7817;
  assign po5767 = new_n7818;
  assign po5768 = new_n7819;
  assign po5769 = new_n7820;
  assign po5770 = new_n7821;
  assign po5771 = new_n7822;
  assign po5772 = new_n7823;
  assign po5773 = new_n7824;
  assign po5774 = new_n7829;
  assign po5775 = new_n7830;
  assign po5776 = new_n7831;
  assign po5777 = new_n7832;
  assign po5778 = new_n7833;
  assign po5779 = new_n7834;
  assign po5780 = new_n7835;
  assign po5781 = new_n7836;
  assign po5782 = new_n7839;
  assign po5783 = new_n7840;
  assign po5784 = new_n7841;
  assign po5785 = new_n7842;
  assign po5786 = new_n7843;
  assign po5787 = new_n7844;
  assign po5788 = new_n7845;
  assign po5789 = new_n7846;
  assign po5790 = new_n7853;
  assign po5791 = new_n7854;
  assign po5792 = new_n7855;
  assign po5793 = new_n7856;
  assign po5794 = new_n7857;
  assign po5795 = new_n7858;
  assign po5796 = new_n7859;
  assign po5797 = new_n7860;
  assign po5798 = new_n7863;
  assign po5799 = new_n7864;
  assign po5800 = new_n7865;
  assign po5801 = new_n7866;
  assign po5802 = new_n7867;
  assign po5803 = new_n7868;
  assign po5804 = new_n7869;
  assign po5805 = new_n7870;
  assign po5806 = new_n7875;
  assign po5807 = new_n7876;
  assign po5808 = new_n7877;
  assign po5809 = new_n7878;
  assign po5810 = new_n7879;
  assign po5811 = new_n7880;
  assign po5812 = new_n7881;
  assign po5813 = new_n7882;
  assign po5814 = new_n7885;
  assign po5815 = new_n7886;
  assign po5816 = new_n7887;
  assign po5817 = new_n7888;
  assign po5818 = new_n7889;
  assign po5819 = new_n7890;
  assign po5820 = new_n7891;
  assign po5821 = new_n7892;
  assign po5822 = new_n7899;
  assign po5823 = new_n7900;
  assign po5824 = new_n7901;
  assign po5825 = new_n7902;
  assign po5826 = new_n7903;
  assign po5827 = new_n7904;
  assign po5828 = new_n7905;
  assign po5829 = new_n7906;
  assign po5830 = new_n7909;
  assign po5831 = new_n7910;
  assign po5832 = new_n7911;
  assign po5833 = new_n7912;
  assign po5834 = new_n7913;
  assign po5835 = new_n7914;
  assign po5836 = new_n7915;
  assign po5837 = new_n7916;
  assign po5838 = new_n7921;
  assign po5839 = new_n7922;
  assign po5840 = new_n7923;
  assign po5841 = new_n7924;
  assign po5842 = new_n7925;
  assign po5843 = new_n7926;
  assign po5844 = new_n7927;
  assign po5845 = new_n7928;
  assign po5846 = new_n7931;
  assign po5847 = new_n7932;
  assign po5848 = new_n7933;
  assign po5849 = new_n7934;
  assign po5850 = new_n7935;
  assign po5851 = new_n7936;
  assign po5852 = new_n7937;
  assign po5853 = new_n7938;
  assign po5854 = new_n7945;
  assign po5855 = new_n7946;
  assign po5856 = new_n7947;
  assign po5857 = new_n7948;
  assign po5858 = new_n7949;
  assign po5859 = new_n7950;
  assign po5860 = new_n7951;
  assign po5861 = new_n7952;
  assign po5862 = new_n7955;
  assign po5863 = new_n7956;
  assign po5864 = new_n7957;
  assign po5865 = new_n7958;
  assign po5866 = new_n7959;
  assign po5867 = new_n7960;
  assign po5868 = new_n7961;
  assign po5869 = new_n7962;
  assign po5870 = new_n7967;
  assign po5871 = new_n7968;
  assign po5872 = new_n7969;
  assign po5873 = new_n7970;
  assign po5874 = new_n7971;
  assign po5875 = new_n7972;
  assign po5876 = new_n7973;
  assign po5877 = new_n7974;
  assign po5878 = new_n7977;
  assign po5879 = new_n7978;
  assign po5880 = new_n7979;
  assign po5881 = new_n7980;
  assign po5882 = new_n7981;
  assign po5883 = new_n7982;
  assign po5884 = new_n7983;
  assign po5885 = new_n7984;
  assign po5886 = new_n7991;
  assign po5887 = new_n7992;
  assign po5888 = new_n7993;
  assign po5889 = new_n7994;
  assign po5890 = new_n7995;
  assign po5891 = new_n7996;
  assign po5892 = new_n7997;
  assign po5893 = new_n7998;
  assign po5894 = new_n8001;
  assign po5895 = new_n8002;
  assign po5896 = new_n8003;
  assign po5897 = new_n8004;
  assign po5898 = new_n8005;
  assign po5899 = new_n8006;
  assign po5900 = new_n8007;
  assign po5901 = new_n8008;
  assign po5902 = new_n8013;
  assign po5903 = new_n8014;
  assign po5904 = new_n8015;
  assign po5905 = new_n8016;
  assign po5906 = new_n8017;
  assign po5907 = new_n8018;
  assign po5908 = new_n8019;
  assign po5909 = new_n8020;
  assign po5910 = new_n8023;
  assign po5911 = new_n8024;
  assign po5912 = new_n8025;
  assign po5913 = new_n8026;
  assign po5914 = new_n8027;
  assign po5915 = new_n8028;
  assign po5916 = new_n8029;
  assign po5917 = new_n8030;
  assign po5918 = new_n8037;
  assign po5919 = new_n8038;
  assign po5920 = new_n8039;
  assign po5921 = new_n8040;
  assign po5922 = new_n8041;
  assign po5923 = new_n8042;
  assign po5924 = new_n8043;
  assign po5925 = new_n8044;
  assign po5926 = new_n8047;
  assign po5927 = new_n8048;
  assign po5928 = new_n8049;
  assign po5929 = new_n8050;
  assign po5930 = new_n8051;
  assign po5931 = new_n8052;
  assign po5932 = new_n8053;
  assign po5933 = new_n8054;
  assign po5934 = new_n8059;
  assign po5935 = new_n8060;
  assign po5936 = new_n8061;
  assign po5937 = new_n8062;
  assign po5938 = new_n8063;
  assign po5939 = new_n8064;
  assign po5940 = new_n8065;
  assign po5941 = new_n8066;
  assign po5942 = new_n8069;
  assign po5943 = new_n8070;
  assign po5944 = new_n8071;
  assign po5945 = new_n8072;
  assign po5946 = new_n8073;
  assign po5947 = new_n8074;
  assign po5948 = new_n8075;
  assign po5949 = new_n8076;
  assign po5950 = new_n8083;
  assign po5951 = new_n8084;
  assign po5952 = new_n8085;
  assign po5953 = new_n8086;
  assign po5954 = new_n8087;
  assign po5955 = new_n8088;
  assign po5956 = new_n8089;
  assign po5957 = new_n8090;
  assign po5958 = new_n8093;
  assign po5959 = new_n8094;
  assign po5960 = new_n8095;
  assign po5961 = new_n8096;
  assign po5962 = new_n8097;
  assign po5963 = new_n8098;
  assign po5964 = new_n8099;
  assign po5965 = new_n8100;
  assign po5966 = new_n8105;
  assign po5967 = new_n8106;
  assign po5968 = new_n8107;
  assign po5969 = new_n8108;
  assign po5970 = new_n8109;
  assign po5971 = new_n8110;
  assign po5972 = new_n8111;
  assign po5973 = new_n8112;
  assign po5974 = new_n8115;
  assign po5975 = new_n8116;
  assign po5976 = new_n8117;
  assign po5977 = new_n8118;
  assign po5978 = new_n8119;
  assign po5979 = new_n8120;
  assign po5980 = new_n8121;
  assign po5981 = new_n8122;
  assign po5982 = new_n8129;
  assign po5983 = new_n8130;
  assign po5984 = new_n8131;
  assign po5985 = new_n8132;
  assign po5986 = new_n8133;
  assign po5987 = new_n8134;
  assign po5988 = new_n8135;
  assign po5989 = new_n8136;
  assign po5990 = new_n8139;
  assign po5991 = new_n8140;
  assign po5992 = new_n8141;
  assign po5993 = new_n8142;
  assign po5994 = new_n8143;
  assign po5995 = new_n8144;
  assign po5996 = new_n8145;
  assign po5997 = new_n8146;
  assign po5998 = new_n8151;
  assign po5999 = new_n8152;
  assign po6000 = new_n8153;
  assign po6001 = new_n8154;
  assign po6002 = new_n8155;
  assign po6003 = new_n8156;
  assign po6004 = new_n8157;
  assign po6005 = new_n8158;
  assign po6006 = new_n8161;
  assign po6007 = new_n8162;
  assign po6008 = new_n8163;
  assign po6009 = new_n8164;
  assign po6010 = new_n8165;
  assign po6011 = new_n8166;
  assign po6012 = new_n8167;
  assign po6013 = new_n8168;
  assign po6014 = new_n8175;
  assign po6015 = new_n8176;
  assign po6016 = new_n8177;
  assign po6017 = new_n8178;
  assign po6018 = new_n8179;
  assign po6019 = new_n8180;
  assign po6020 = new_n8181;
  assign po6021 = new_n8182;
  assign po6022 = new_n8185;
  assign po6023 = new_n8186;
  assign po6024 = new_n8187;
  assign po6025 = new_n8188;
  assign po6026 = new_n8189;
  assign po6027 = new_n8190;
  assign po6028 = new_n8191;
  assign po6029 = new_n8192;
  assign po6030 = new_n8197;
  assign po6031 = new_n8198;
  assign po6032 = new_n8199;
  assign po6033 = new_n8200;
  assign po6034 = new_n8201;
  assign po6035 = new_n8202;
  assign po6036 = new_n8203;
  assign po6037 = new_n8204;
  assign po6038 = new_n8207;
  assign po6039 = new_n8208;
  assign po6040 = new_n8209;
  assign po6041 = new_n8210;
  assign po6042 = new_n8211;
  assign po6043 = new_n8212;
  assign po6044 = new_n8213;
  assign po6045 = new_n8214;
  assign po6046 = new_n8221;
  assign po6047 = new_n8222;
  assign po6048 = new_n8223;
  assign po6049 = new_n8224;
  assign po6050 = new_n8225;
  assign po6051 = new_n8226;
  assign po6052 = new_n8227;
  assign po6053 = new_n8228;
  assign po6054 = new_n8231;
  assign po6055 = new_n8232;
  assign po6056 = new_n8233;
  assign po6057 = new_n8234;
  assign po6058 = new_n8235;
  assign po6059 = new_n8236;
  assign po6060 = new_n8237;
  assign po6061 = new_n8238;
  assign po6062 = new_n8243;
  assign po6063 = new_n8244;
  assign po6064 = new_n8245;
  assign po6065 = new_n8246;
  assign po6066 = new_n8247;
  assign po6067 = new_n8248;
  assign po6068 = new_n8249;
  assign po6069 = new_n8250;
  assign po6070 = new_n8253;
  assign po6071 = new_n8254;
  assign po6072 = new_n8255;
  assign po6073 = new_n8256;
  assign po6074 = new_n8257;
  assign po6075 = new_n8258;
  assign po6076 = new_n8259;
  assign po6077 = new_n8260;
  assign po6078 = new_n8267;
  assign po6079 = new_n8268;
  assign po6080 = new_n8269;
  assign po6081 = new_n8270;
  assign po6082 = new_n8271;
  assign po6083 = new_n8272;
  assign po6084 = new_n8273;
  assign po6085 = new_n8274;
  assign po6086 = new_n8277;
  assign po6087 = new_n8278;
  assign po6088 = new_n8279;
  assign po6089 = new_n8280;
  assign po6090 = new_n8281;
  assign po6091 = new_n8282;
  assign po6092 = new_n8283;
  assign po6093 = new_n8284;
  assign po6094 = new_n8289;
  assign po6095 = new_n8290;
  assign po6096 = new_n8291;
  assign po6097 = new_n8292;
  assign po6098 = new_n8293;
  assign po6099 = new_n8294;
  assign po6100 = new_n8295;
  assign po6101 = new_n8296;
  assign po6102 = new_n8299;
  assign po6103 = new_n8300;
  assign po6104 = new_n8301;
  assign po6105 = new_n8302;
  assign po6106 = new_n8303;
  assign po6107 = new_n8304;
  assign po6108 = new_n8305;
  assign po6109 = new_n8306;
  assign po6110 = new_n8313;
  assign po6111 = new_n8314;
  assign po6112 = new_n8315;
  assign po6113 = new_n8316;
  assign po6114 = new_n8317;
  assign po6115 = new_n8318;
  assign po6116 = new_n8319;
  assign po6117 = new_n8320;
  assign po6118 = new_n8323;
  assign po6119 = new_n8324;
  assign po6120 = new_n8325;
  assign po6121 = new_n8326;
  assign po6122 = new_n8327;
  assign po6123 = new_n8328;
  assign po6124 = new_n8329;
  assign po6125 = new_n8330;
  assign po6126 = new_n8335;
  assign po6127 = new_n8336;
  assign po6128 = new_n8337;
  assign po6129 = new_n8338;
  assign po6130 = new_n8339;
  assign po6131 = new_n8340;
  assign po6132 = new_n8341;
  assign po6133 = new_n8342;
  assign po6134 = new_n8345;
  assign po6135 = new_n8346;
  assign po6136 = new_n8347;
  assign po6137 = new_n8348;
  assign po6138 = new_n8349;
  assign po6139 = new_n8350;
  assign po6140 = new_n8351;
  assign po6141 = new_n8352;
  assign po6142 = new_n8359;
  assign po6143 = new_n8360;
  assign po6144 = new_n8361;
  assign po6145 = new_n8362;
  assign po6146 = new_n8363;
  assign po6147 = new_n8364;
  assign po6148 = new_n8365;
  assign po6149 = new_n8366;
  assign po6150 = new_n8369;
  assign po6151 = new_n8370;
  assign po6152 = new_n8371;
  assign po6153 = new_n8372;
  assign po6154 = new_n8373;
  assign po6155 = new_n8374;
  assign po6156 = new_n8375;
  assign po6157 = new_n8376;
  assign po6158 = new_n8381;
  assign po6159 = new_n8382;
  assign po6160 = new_n8383;
  assign po6161 = new_n8384;
  assign po6162 = new_n8385;
  assign po6163 = new_n8386;
  assign po6164 = new_n8387;
  assign po6165 = new_n8388;
  assign po6166 = new_n8391;
  assign po6167 = new_n8392;
  assign po6168 = new_n8393;
  assign po6169 = new_n8394;
  assign po6170 = new_n8395;
  assign po6171 = new_n8396;
  assign po6172 = new_n8397;
  assign po6173 = new_n8398;
  assign po6174 = new_n9311;
  assign po6175 = new_n10089;
  assign po6176 = new_n10871;
  assign po6177 = new_n11649;
  assign po6178 = new_n12427;
  assign po6179 = new_n13205;
  assign po6180 = new_n13983;
  assign po6181 = new_n14761;
  assign po6182 = new_n14772;
  assign po6183 = new_n14782;
  assign po6184 = new_n14792;
  assign po6185 = new_n14802;
  assign po6186 = new_n14812;
  assign po6187 = new_n14822;
  assign po6188 = new_n14832;
  assign po6189 = new_n14842;
  assign po6190 = new_n14852;
  assign po6191 = new_n14859;
  assign po6192 = new_n14866;
  assign po6193 = new_n14873;
  assign po6194 = new_n14880;
  assign po6195 = new_n14887;
  assign po6196 = new_n14894;
  assign po6197 = new_n14901;
  assign po6198 = new_n14908;
  assign po6199 = new_n14915;
  assign po6200 = new_n14922;
  assign po6201 = new_n14929;
  assign po6202 = new_n14936;
  assign po6203 = new_n14943;
  assign po6204 = new_n14950;
  assign po6205 = new_n14957;
  assign po6206 = new_n14961;
  assign po6207 = new_n14962;
  assign po6208 = new_n14963;
  assign po6209 = new_n14964;
  assign po6210 = new_n14965;
  assign po6211 = new_n14966;
  assign po6212 = new_n14967;
  assign po6213 = new_n14968;
  assign po6214 = new_n14969;
  assign po6215 = new_n14970;
  assign po6216 = new_n14971;
  assign po6217 = new_n14972;
  assign po6218 = new_n14973;
  assign po6219 = new_n14974;
  assign po6220 = new_n14975;
  assign po6221 = new_n14976;
  assign po6222 = new_n14977;
  assign po6223 = new_n14978;
  assign po6224 = new_n14979;
  assign po6225 = new_n14980;
  assign po6226 = new_n14981;
  assign po6227 = new_n14982;
  assign po6228 = new_n14983;
  assign po6229 = new_n14984;
  assign po6230 = new_n14985;
  assign po6231 = new_n14986;
  assign po6232 = new_n14987;
  assign po6233 = new_n14988;
  assign po6234 = new_n14989;
  assign po6235 = new_n14990;
  assign po6236 = new_n14991;
  assign po6237 = new_n14992;
  assign po6238 = new_n14996;
  assign po6239 = new_n14997;
  assign po6240 = new_n14998;
  assign po6241 = new_n14999;
  assign po6242 = new_n15000;
  assign po6243 = new_n15001;
  assign po6244 = new_n15002;
  assign po6245 = new_n15003;
  assign po6246 = new_n15004;
  assign po6247 = new_n15005;
  assign po6248 = new_n15006;
  assign po6249 = new_n15007;
  assign po6250 = new_n15008;
  assign po6251 = new_n15009;
  assign po6252 = new_n15010;
  assign po6253 = new_n15011;
  assign po6254 = new_n15012;
  assign po6255 = new_n15013;
  assign po6256 = new_n15014;
  assign po6257 = new_n15015;
  assign po6258 = new_n15016;
  assign po6259 = new_n15017;
  assign po6260 = new_n15018;
  assign po6261 = new_n15019;
  assign po6262 = new_n15020;
  assign po6263 = new_n15021;
  assign po6264 = new_n15022;
  assign po6265 = new_n15023;
  assign po6266 = new_n15024;
  assign po6267 = new_n15025;
  assign po6268 = new_n15026;
  assign po6269 = new_n15027;
  assign po6270 = new_n15031;
  assign po6271 = new_n15032;
  assign po6272 = new_n15033;
  assign po6273 = new_n15034;
  assign po6274 = new_n15035;
  assign po6275 = new_n15036;
  assign po6276 = new_n15037;
  assign po6277 = new_n15038;
  assign po6278 = new_n15039;
  assign po6279 = new_n15040;
  assign po6280 = new_n15041;
  assign po6281 = new_n15042;
  assign po6282 = new_n15043;
  assign po6283 = new_n15044;
  assign po6284 = new_n15045;
  assign po6285 = new_n15046;
  assign po6286 = new_n15047;
  assign po6287 = new_n15048;
  assign po6288 = new_n15049;
  assign po6289 = new_n15050;
  assign po6290 = new_n15051;
  assign po6291 = new_n15052;
  assign po6292 = new_n15053;
  assign po6293 = new_n15054;
  assign po6294 = new_n15055;
  assign po6295 = new_n15056;
  assign po6296 = new_n15057;
  assign po6297 = new_n15058;
  assign po6298 = new_n15059;
  assign po6299 = new_n15060;
  assign po6300 = new_n15061;
  assign po6301 = new_n15062;
  assign po6302 = new_n15064;
  assign po6303 = new_n15065;
  assign po6304 = new_n15066;
  assign po6305 = new_n15067;
  assign po6306 = new_n15068;
  assign po6307 = new_n15069;
  assign po6308 = new_n15070;
  assign po6309 = new_n15071;
  assign po6310 = new_n15072;
  assign po6311 = new_n15073;
  assign po6312 = new_n15074;
  assign po6313 = new_n15075;
  assign po6314 = new_n15076;
  assign po6315 = new_n15077;
  assign po6316 = new_n15078;
  assign po6317 = new_n15079;
  assign po6318 = new_n15080;
  assign po6319 = new_n15081;
  assign po6320 = new_n15082;
  assign po6321 = new_n15083;
  assign po6322 = new_n15084;
  assign po6323 = new_n15085;
  assign po6324 = new_n15086;
  assign po6325 = new_n15087;
  assign po6326 = new_n15088;
  assign po6327 = new_n15089;
  assign po6328 = new_n15090;
  assign po6329 = new_n15091;
  assign po6330 = new_n15092;
  assign po6331 = new_n15093;
  assign po6332 = new_n15094;
  assign po6333 = new_n15095;
  assign po6334 = new_n15097;
  assign po6335 = new_n15098;
  assign po6336 = new_n15099;
  assign po6337 = new_n15100;
  assign po6338 = new_n15101;
  assign po6339 = new_n15102;
  assign po6340 = new_n15103;
  assign po6341 = new_n15104;
  assign po6342 = new_n15105;
  assign po6343 = new_n15106;
  assign po6344 = new_n15107;
  assign po6345 = new_n15108;
  assign po6346 = new_n15109;
  assign po6347 = new_n15110;
  assign po6348 = new_n15111;
  assign po6349 = new_n15112;
  assign po6350 = new_n15113;
  assign po6351 = new_n15114;
  assign po6352 = new_n15115;
  assign po6353 = new_n15116;
  assign po6354 = new_n15117;
  assign po6355 = new_n15118;
  assign po6356 = new_n15119;
  assign po6357 = new_n15120;
  assign po6358 = new_n15121;
  assign po6359 = new_n15122;
  assign po6360 = new_n15123;
  assign po6361 = new_n15124;
  assign po6362 = new_n15125;
  assign po6363 = new_n15126;
  assign po6364 = new_n15127;
  assign po6365 = new_n15128;
  assign po6366 = new_n15130;
  assign po6367 = new_n15131;
  assign po6368 = new_n15132;
  assign po6369 = new_n15133;
  assign po6370 = new_n15134;
  assign po6371 = new_n15135;
  assign po6372 = new_n15136;
  assign po6373 = new_n15137;
  assign po6374 = new_n15138;
  assign po6375 = new_n15139;
  assign po6376 = new_n15140;
  assign po6377 = new_n15141;
  assign po6378 = new_n15142;
  assign po6379 = new_n15143;
  assign po6380 = new_n15144;
  assign po6381 = new_n15145;
  assign po6382 = new_n15146;
  assign po6383 = new_n15147;
  assign po6384 = new_n15148;
  assign po6385 = new_n15149;
  assign po6386 = new_n15150;
  assign po6387 = new_n15151;
  assign po6388 = new_n15152;
  assign po6389 = new_n15153;
  assign po6390 = new_n15154;
  assign po6391 = new_n15155;
  assign po6392 = new_n15156;
  assign po6393 = new_n15157;
  assign po6394 = new_n15158;
  assign po6395 = new_n15159;
  assign po6396 = new_n15160;
  assign po6397 = new_n15161;
  assign po6398 = new_n15164;
  assign po6399 = new_n15165;
  assign po6400 = new_n15166;
  assign po6401 = new_n15167;
  assign po6402 = new_n15168;
  assign po6403 = new_n15169;
  assign po6404 = new_n15170;
  assign po6405 = new_n15171;
  assign po6406 = new_n15172;
  assign po6407 = new_n15173;
  assign po6408 = new_n15174;
  assign po6409 = new_n15175;
  assign po6410 = new_n15176;
  assign po6411 = new_n15177;
  assign po6412 = new_n15178;
  assign po6413 = new_n15179;
  assign po6414 = new_n15180;
  assign po6415 = new_n15181;
  assign po6416 = new_n15182;
  assign po6417 = new_n15183;
  assign po6418 = new_n15184;
  assign po6419 = new_n15185;
  assign po6420 = new_n15186;
  assign po6421 = new_n15187;
  assign po6422 = new_n15188;
  assign po6423 = new_n15189;
  assign po6424 = new_n15190;
  assign po6425 = new_n15191;
  assign po6426 = new_n15192;
  assign po6427 = new_n15193;
  assign po6428 = new_n15194;
  assign po6429 = new_n15195;
  assign po6430 = new_n15197;
  assign po6431 = new_n15198;
  assign po6432 = new_n15199;
  assign po6433 = new_n15200;
  assign po6434 = new_n15201;
  assign po6435 = new_n15202;
  assign po6436 = new_n15203;
  assign po6437 = new_n15204;
  assign po6438 = new_n15205;
  assign po6439 = new_n15206;
  assign po6440 = new_n15207;
  assign po6441 = new_n15208;
  assign po6442 = new_n15209;
  assign po6443 = new_n15210;
  assign po6444 = new_n15211;
  assign po6445 = new_n15212;
  assign po6446 = new_n15213;
  assign po6447 = new_n15214;
  assign po6448 = new_n15215;
  assign po6449 = new_n15216;
  assign po6450 = new_n15217;
  assign po6451 = new_n15218;
  assign po6452 = new_n15219;
  assign po6453 = new_n15220;
  assign po6454 = new_n15221;
  assign po6455 = new_n15222;
  assign po6456 = new_n15223;
  assign po6457 = new_n15224;
  assign po6458 = new_n15225;
  assign po6459 = new_n15226;
  assign po6460 = new_n15227;
  assign po6461 = new_n15228;
  assign po6462 = new_n15230;
  assign po6463 = new_n15231;
  assign po6464 = new_n15232;
  assign po6465 = new_n15233;
  assign po6466 = new_n15234;
  assign po6467 = new_n15235;
  assign po6468 = new_n15236;
  assign po6469 = new_n15237;
  assign po6470 = new_n15238;
  assign po6471 = new_n15239;
  assign po6472 = new_n15240;
  assign po6473 = new_n15241;
  assign po6474 = new_n15242;
  assign po6475 = new_n15243;
  assign po6476 = new_n15244;
  assign po6477 = new_n15245;
  assign po6478 = new_n15246;
  assign po6479 = new_n15247;
  assign po6480 = new_n15248;
  assign po6481 = new_n15249;
  assign po6482 = new_n15250;
  assign po6483 = new_n15251;
  assign po6484 = new_n15252;
  assign po6485 = new_n15253;
  assign po6486 = new_n15254;
  assign po6487 = new_n15255;
  assign po6488 = new_n15256;
  assign po6489 = new_n15257;
  assign po6490 = new_n15258;
  assign po6491 = new_n15259;
  assign po6492 = new_n15260;
  assign po6493 = new_n15261;
  assign po6494 = new_n15263;
  assign po6495 = new_n15264;
  assign po6496 = new_n15265;
  assign po6497 = new_n15266;
  assign po6498 = new_n15267;
  assign po6499 = new_n15268;
  assign po6500 = new_n15269;
  assign po6501 = new_n15270;
  assign po6502 = new_n15271;
  assign po6503 = new_n15272;
  assign po6504 = new_n15273;
  assign po6505 = new_n15274;
  assign po6506 = new_n15275;
  assign po6507 = new_n15276;
  assign po6508 = new_n15277;
  assign po6509 = new_n15278;
  assign po6510 = new_n15279;
  assign po6511 = new_n15280;
  assign po6512 = new_n15281;
  assign po6513 = new_n15282;
  assign po6514 = new_n15283;
  assign po6515 = new_n15284;
  assign po6516 = new_n15285;
  assign po6517 = new_n15286;
  assign po6518 = new_n15287;
  assign po6519 = new_n15288;
  assign po6520 = new_n15289;
  assign po6521 = new_n15290;
  assign po6522 = new_n15291;
  assign po6523 = new_n15292;
  assign po6524 = new_n15293;
  assign po6525 = new_n15294;
  assign po6526 = new_n15296;
  assign po6527 = new_n15297;
  assign po6528 = new_n15298;
  assign po6529 = new_n15299;
  assign po6530 = new_n15300;
  assign po6531 = new_n15301;
  assign po6532 = new_n15302;
  assign po6533 = new_n15303;
  assign po6534 = new_n15304;
  assign po6535 = new_n15305;
  assign po6536 = new_n15306;
  assign po6537 = new_n15307;
  assign po6538 = new_n15308;
  assign po6539 = new_n15309;
  assign po6540 = new_n15310;
  assign po6541 = new_n15311;
  assign po6542 = new_n15312;
  assign po6543 = new_n15313;
  assign po6544 = new_n15314;
  assign po6545 = new_n15315;
  assign po6546 = new_n15316;
  assign po6547 = new_n15317;
  assign po6548 = new_n15318;
  assign po6549 = new_n15319;
  assign po6550 = new_n15320;
  assign po6551 = new_n15321;
  assign po6552 = new_n15322;
  assign po6553 = new_n15323;
  assign po6554 = new_n15324;
  assign po6555 = new_n15325;
  assign po6556 = new_n15326;
  assign po6557 = new_n15327;
  assign po6558 = new_n15329;
  assign po6559 = new_n15330;
  assign po6560 = new_n15331;
  assign po6561 = new_n15332;
  assign po6562 = new_n15333;
  assign po6563 = new_n15334;
  assign po6564 = new_n15335;
  assign po6565 = new_n15336;
  assign po6566 = new_n15337;
  assign po6567 = new_n15338;
  assign po6568 = new_n15339;
  assign po6569 = new_n15340;
  assign po6570 = new_n15341;
  assign po6571 = new_n15342;
  assign po6572 = new_n15343;
  assign po6573 = new_n15344;
  assign po6574 = new_n15345;
  assign po6575 = new_n15346;
  assign po6576 = new_n15347;
  assign po6577 = new_n15348;
  assign po6578 = new_n15349;
  assign po6579 = new_n15350;
  assign po6580 = new_n15351;
  assign po6581 = new_n15352;
  assign po6582 = new_n15353;
  assign po6583 = new_n15354;
  assign po6584 = new_n15355;
  assign po6585 = new_n15356;
  assign po6586 = new_n15357;
  assign po6587 = new_n15358;
  assign po6588 = new_n15359;
  assign po6589 = new_n15360;
  assign po6590 = new_n15362;
  assign po6591 = new_n15363;
  assign po6592 = new_n15364;
  assign po6593 = new_n15365;
  assign po6594 = new_n15366;
  assign po6595 = new_n15367;
  assign po6596 = new_n15368;
  assign po6597 = new_n15369;
  assign po6598 = new_n15370;
  assign po6599 = new_n15371;
  assign po6600 = new_n15372;
  assign po6601 = new_n15373;
  assign po6602 = new_n15374;
  assign po6603 = new_n15375;
  assign po6604 = new_n15376;
  assign po6605 = new_n15377;
  assign po6606 = new_n15378;
  assign po6607 = new_n15379;
  assign po6608 = new_n15380;
  assign po6609 = new_n15381;
  assign po6610 = new_n15382;
  assign po6611 = new_n15383;
  assign po6612 = new_n15384;
  assign po6613 = new_n15385;
  assign po6614 = new_n15386;
  assign po6615 = new_n15387;
  assign po6616 = new_n15388;
  assign po6617 = new_n15389;
  assign po6618 = new_n15390;
  assign po6619 = new_n15391;
  assign po6620 = new_n15392;
  assign po6621 = new_n15393;
  assign po6622 = new_n15395;
  assign po6623 = new_n15396;
  assign po6624 = new_n15397;
  assign po6625 = new_n15398;
  assign po6626 = new_n15399;
  assign po6627 = new_n15400;
  assign po6628 = new_n15401;
  assign po6629 = new_n15402;
  assign po6630 = new_n15403;
  assign po6631 = new_n15404;
  assign po6632 = new_n15405;
  assign po6633 = new_n15406;
  assign po6634 = new_n15407;
  assign po6635 = new_n15408;
  assign po6636 = new_n15409;
  assign po6637 = new_n15410;
  assign po6638 = new_n15411;
  assign po6639 = new_n15412;
  assign po6640 = new_n15413;
  assign po6641 = new_n15414;
  assign po6642 = new_n15415;
  assign po6643 = new_n15416;
  assign po6644 = new_n15417;
  assign po6645 = new_n15418;
  assign po6646 = new_n15419;
  assign po6647 = new_n15420;
  assign po6648 = new_n15421;
  assign po6649 = new_n15422;
  assign po6650 = new_n15423;
  assign po6651 = new_n15424;
  assign po6652 = new_n15425;
  assign po6653 = new_n15426;
  assign po6654 = new_n15428;
  assign po6655 = new_n15429;
  assign po6656 = new_n15430;
  assign po6657 = new_n15431;
  assign po6658 = new_n15432;
  assign po6659 = new_n15433;
  assign po6660 = new_n15434;
  assign po6661 = new_n15435;
  assign po6662 = new_n15436;
  assign po6663 = new_n15437;
  assign po6664 = new_n15438;
  assign po6665 = new_n15439;
  assign po6666 = new_n15440;
  assign po6667 = new_n15441;
  assign po6668 = new_n15442;
  assign po6669 = new_n15443;
  assign po6670 = new_n15444;
  assign po6671 = new_n15445;
  assign po6672 = new_n15446;
  assign po6673 = new_n15447;
  assign po6674 = new_n15448;
  assign po6675 = new_n15449;
  assign po6676 = new_n15450;
  assign po6677 = new_n15451;
  assign po6678 = new_n15452;
  assign po6679 = new_n15453;
  assign po6680 = new_n15454;
  assign po6681 = new_n15455;
  assign po6682 = new_n15456;
  assign po6683 = new_n15457;
  assign po6684 = new_n15458;
  assign po6685 = new_n15459;
  assign po6686 = new_n15461;
  assign po6687 = new_n15462;
  assign po6688 = new_n15463;
  assign po6689 = new_n15464;
  assign po6690 = new_n15465;
  assign po6691 = new_n15466;
  assign po6692 = new_n15467;
  assign po6693 = new_n15468;
  assign po6694 = new_n15469;
  assign po6695 = new_n15470;
  assign po6696 = new_n15471;
  assign po6697 = new_n15472;
  assign po6698 = new_n15473;
  assign po6699 = new_n15474;
  assign po6700 = new_n15475;
  assign po6701 = new_n15476;
  assign po6702 = new_n15477;
  assign po6703 = new_n15478;
  assign po6704 = new_n15479;
  assign po6705 = new_n15480;
  assign po6706 = new_n15481;
  assign po6707 = new_n15482;
  assign po6708 = new_n15483;
  assign po6709 = new_n15484;
  assign po6710 = new_n15485;
  assign po6711 = new_n15486;
  assign po6712 = new_n15487;
  assign po6713 = new_n15488;
  assign po6714 = new_n15489;
  assign po6715 = new_n15490;
  assign po6716 = new_n15491;
  assign po6717 = new_n15492;
  assign po6718 = new_n15494;
  assign po6719 = new_n15495;
  assign po6720 = new_n15496;
  assign po6721 = new_n15497;
  assign po6722 = new_n15498;
  assign po6723 = new_n15499;
  assign po6724 = new_n15500;
  assign po6725 = new_n15501;
  assign po6726 = new_n15502;
  assign po6727 = new_n15503;
  assign po6728 = new_n15504;
  assign po6729 = new_n15505;
  assign po6730 = new_n15506;
  assign po6731 = new_n15507;
  assign po6732 = new_n15508;
  assign po6733 = new_n15509;
  assign po6734 = new_n15510;
  assign po6735 = new_n15511;
  assign po6736 = new_n15512;
  assign po6737 = new_n15513;
  assign po6738 = new_n15514;
  assign po6739 = new_n15515;
  assign po6740 = new_n15516;
  assign po6741 = new_n15517;
  assign po6742 = new_n15518;
  assign po6743 = new_n15519;
  assign po6744 = new_n15520;
  assign po6745 = new_n15521;
  assign po6746 = new_n15522;
  assign po6747 = new_n15523;
  assign po6748 = new_n15524;
  assign po6749 = new_n15525;
  assign po6750 = new_n15527;
  assign po6751 = new_n15528;
  assign po6752 = new_n15529;
  assign po6753 = new_n15530;
  assign po6754 = new_n15531;
  assign po6755 = new_n15532;
  assign po6756 = new_n15533;
  assign po6757 = new_n15534;
  assign po6758 = new_n15535;
  assign po6759 = new_n15536;
  assign po6760 = new_n15537;
  assign po6761 = new_n15538;
  assign po6762 = new_n15539;
  assign po6763 = new_n15540;
  assign po6764 = new_n15541;
  assign po6765 = new_n15542;
  assign po6766 = new_n15543;
  assign po6767 = new_n15544;
  assign po6768 = new_n15545;
  assign po6769 = new_n15546;
  assign po6770 = new_n15547;
  assign po6771 = new_n15548;
  assign po6772 = new_n15549;
  assign po6773 = new_n15550;
  assign po6774 = new_n15551;
  assign po6775 = new_n15552;
  assign po6776 = new_n15553;
  assign po6777 = new_n15554;
  assign po6778 = new_n15555;
  assign po6779 = new_n15556;
  assign po6780 = new_n15557;
  assign po6781 = new_n15558;
  assign po6782 = new_n15560;
  assign po6783 = new_n15561;
  assign po6784 = new_n15562;
  assign po6785 = new_n15563;
  assign po6786 = new_n15564;
  assign po6787 = new_n15565;
  assign po6788 = new_n15566;
  assign po6789 = new_n15567;
  assign po6790 = new_n15568;
  assign po6791 = new_n15569;
  assign po6792 = new_n15570;
  assign po6793 = new_n15571;
  assign po6794 = new_n15572;
  assign po6795 = new_n15573;
  assign po6796 = new_n15574;
  assign po6797 = new_n15575;
  assign po6798 = new_n15576;
  assign po6799 = new_n15577;
  assign po6800 = new_n15578;
  assign po6801 = new_n15579;
  assign po6802 = new_n15580;
  assign po6803 = new_n15581;
  assign po6804 = new_n15582;
  assign po6805 = new_n15583;
  assign po6806 = new_n15584;
  assign po6807 = new_n15585;
  assign po6808 = new_n15586;
  assign po6809 = new_n15587;
  assign po6810 = new_n15588;
  assign po6811 = new_n15589;
  assign po6812 = new_n15590;
  assign po6813 = new_n15591;
  assign po6814 = new_n15593;
  assign po6815 = new_n15594;
  assign po6816 = new_n15595;
  assign po6817 = new_n15596;
  assign po6818 = new_n15597;
  assign po6819 = new_n15598;
  assign po6820 = new_n15599;
  assign po6821 = new_n15600;
  assign po6822 = new_n15601;
  assign po6823 = new_n15602;
  assign po6824 = new_n15603;
  assign po6825 = new_n15604;
  assign po6826 = new_n15605;
  assign po6827 = new_n15606;
  assign po6828 = new_n15607;
  assign po6829 = new_n15608;
  assign po6830 = new_n15609;
  assign po6831 = new_n15610;
  assign po6832 = new_n15611;
  assign po6833 = new_n15612;
  assign po6834 = new_n15613;
  assign po6835 = new_n15614;
  assign po6836 = new_n15615;
  assign po6837 = new_n15616;
  assign po6838 = new_n15617;
  assign po6839 = new_n15618;
  assign po6840 = new_n15619;
  assign po6841 = new_n15620;
  assign po6842 = new_n15621;
  assign po6843 = new_n15622;
  assign po6844 = new_n15623;
  assign po6845 = new_n15624;
  assign po6846 = new_n15626;
  assign po6847 = new_n15627;
  assign po6848 = new_n15628;
  assign po6849 = new_n15629;
  assign po6850 = new_n15630;
  assign po6851 = new_n15631;
  assign po6852 = new_n15632;
  assign po6853 = new_n15633;
  assign po6854 = new_n15634;
  assign po6855 = new_n15635;
  assign po6856 = new_n15636;
  assign po6857 = new_n15637;
  assign po6858 = new_n15638;
  assign po6859 = new_n15639;
  assign po6860 = new_n15640;
  assign po6861 = new_n15641;
  assign po6862 = new_n15642;
  assign po6863 = new_n15643;
  assign po6864 = new_n15644;
  assign po6865 = new_n15645;
  assign po6866 = new_n15646;
  assign po6867 = new_n15647;
  assign po6868 = new_n15648;
  assign po6869 = new_n15649;
  assign po6870 = new_n15650;
  assign po6871 = new_n15651;
  assign po6872 = new_n15652;
  assign po6873 = new_n15653;
  assign po6874 = new_n15654;
  assign po6875 = new_n15655;
  assign po6876 = new_n15656;
  assign po6877 = new_n15657;
  assign po6878 = new_n15659;
  assign po6879 = new_n15660;
  assign po6880 = new_n15661;
  assign po6881 = new_n15662;
  assign po6882 = new_n15663;
  assign po6883 = new_n15664;
  assign po6884 = new_n15665;
  assign po6885 = new_n15666;
  assign po6886 = new_n15667;
  assign po6887 = new_n15668;
  assign po6888 = new_n15669;
  assign po6889 = new_n15670;
  assign po6890 = new_n15671;
  assign po6891 = new_n15672;
  assign po6892 = new_n15673;
  assign po6893 = new_n15674;
  assign po6894 = new_n15675;
  assign po6895 = new_n15676;
  assign po6896 = new_n15677;
  assign po6897 = new_n15678;
  assign po6898 = new_n15679;
  assign po6899 = new_n15680;
  assign po6900 = new_n15681;
  assign po6901 = new_n15682;
  assign po6902 = new_n15683;
  assign po6903 = new_n15684;
  assign po6904 = new_n15685;
  assign po6905 = new_n15686;
  assign po6906 = new_n15687;
  assign po6907 = new_n15688;
  assign po6908 = new_n15689;
  assign po6909 = new_n15690;
  assign po6910 = new_n15692;
  assign po6911 = new_n15693;
  assign po6912 = new_n15694;
  assign po6913 = new_n15695;
  assign po6914 = new_n15696;
  assign po6915 = new_n15697;
  assign po6916 = new_n15698;
  assign po6917 = new_n15699;
  assign po6918 = new_n15700;
  assign po6919 = new_n15701;
  assign po6920 = new_n15702;
  assign po6921 = new_n15703;
  assign po6922 = new_n15704;
  assign po6923 = new_n15705;
  assign po6924 = new_n15706;
  assign po6925 = new_n15707;
  assign po6926 = new_n15708;
  assign po6927 = new_n15709;
  assign po6928 = new_n15710;
  assign po6929 = new_n15711;
  assign po6930 = new_n15712;
  assign po6931 = new_n15713;
  assign po6932 = new_n15714;
  assign po6933 = new_n15715;
  assign po6934 = new_n15716;
  assign po6935 = new_n15717;
  assign po6936 = new_n15718;
  assign po6937 = new_n15719;
  assign po6938 = new_n15720;
  assign po6939 = new_n15721;
  assign po6940 = new_n15722;
  assign po6941 = new_n15723;
  assign po6942 = new_n15725;
  assign po6943 = new_n15726;
  assign po6944 = new_n15727;
  assign po6945 = new_n15728;
  assign po6946 = new_n15729;
  assign po6947 = new_n15730;
  assign po6948 = new_n15731;
  assign po6949 = new_n15732;
  assign po6950 = new_n15733;
  assign po6951 = new_n15734;
  assign po6952 = new_n15735;
  assign po6953 = new_n15736;
  assign po6954 = new_n15737;
  assign po6955 = new_n15738;
  assign po6956 = new_n15739;
  assign po6957 = new_n15740;
  assign po6958 = new_n15741;
  assign po6959 = new_n15742;
  assign po6960 = new_n15743;
  assign po6961 = new_n15744;
  assign po6962 = new_n15745;
  assign po6963 = new_n15746;
  assign po6964 = new_n15747;
  assign po6965 = new_n15748;
  assign po6966 = new_n15749;
  assign po6967 = new_n15750;
  assign po6968 = new_n15751;
  assign po6969 = new_n15752;
  assign po6970 = new_n15753;
  assign po6971 = new_n15754;
  assign po6972 = new_n15755;
  assign po6973 = new_n15756;
  assign po6974 = new_n15758;
  assign po6975 = new_n15759;
  assign po6976 = new_n15760;
  assign po6977 = new_n15761;
  assign po6978 = new_n15762;
  assign po6979 = new_n15763;
  assign po6980 = new_n15764;
  assign po6981 = new_n15765;
  assign po6982 = new_n15766;
  assign po6983 = new_n15767;
  assign po6984 = new_n15768;
  assign po6985 = new_n15769;
  assign po6986 = new_n15770;
  assign po6987 = new_n15771;
  assign po6988 = new_n15772;
  assign po6989 = new_n15773;
  assign po6990 = new_n15774;
  assign po6991 = new_n15775;
  assign po6992 = new_n15776;
  assign po6993 = new_n15777;
  assign po6994 = new_n15778;
  assign po6995 = new_n15779;
  assign po6996 = new_n15780;
  assign po6997 = new_n15781;
  assign po6998 = new_n15782;
  assign po6999 = new_n15783;
  assign po7000 = new_n15784;
  assign po7001 = new_n15785;
  assign po7002 = new_n15786;
  assign po7003 = new_n15787;
  assign po7004 = new_n15788;
  assign po7005 = new_n15789;
  assign po7006 = new_n15791;
  assign po7007 = new_n15792;
  assign po7008 = new_n15793;
  assign po7009 = new_n15794;
  assign po7010 = new_n15795;
  assign po7011 = new_n15796;
  assign po7012 = new_n15797;
  assign po7013 = new_n15798;
  assign po7014 = new_n15799;
  assign po7015 = new_n15800;
  assign po7016 = new_n15801;
  assign po7017 = new_n15802;
  assign po7018 = new_n15803;
  assign po7019 = new_n15804;
  assign po7020 = new_n15805;
  assign po7021 = new_n15806;
  assign po7022 = new_n15807;
  assign po7023 = new_n15808;
  assign po7024 = new_n15809;
  assign po7025 = new_n15810;
  assign po7026 = new_n15811;
  assign po7027 = new_n15812;
  assign po7028 = new_n15813;
  assign po7029 = new_n15814;
  assign po7030 = new_n15815;
  assign po7031 = new_n15816;
  assign po7032 = new_n15817;
  assign po7033 = new_n15818;
  assign po7034 = new_n15819;
  assign po7035 = new_n15820;
  assign po7036 = new_n15821;
  assign po7037 = new_n15822;
  assign po7038 = new_n15824;
  assign po7039 = new_n15825;
  assign po7040 = new_n15826;
  assign po7041 = new_n15827;
  assign po7042 = new_n15828;
  assign po7043 = new_n15829;
  assign po7044 = new_n15830;
  assign po7045 = new_n15831;
  assign po7046 = new_n15832;
  assign po7047 = new_n15833;
  assign po7048 = new_n15834;
  assign po7049 = new_n15835;
  assign po7050 = new_n15836;
  assign po7051 = new_n15837;
  assign po7052 = new_n15838;
  assign po7053 = new_n15839;
  assign po7054 = new_n15840;
  assign po7055 = new_n15841;
  assign po7056 = new_n15842;
  assign po7057 = new_n15843;
  assign po7058 = new_n15844;
  assign po7059 = new_n15845;
  assign po7060 = new_n15846;
  assign po7061 = new_n15847;
  assign po7062 = new_n15848;
  assign po7063 = new_n15849;
  assign po7064 = new_n15850;
  assign po7065 = new_n15851;
  assign po7066 = new_n15852;
  assign po7067 = new_n15853;
  assign po7068 = new_n15854;
  assign po7069 = new_n15855;
  assign po7070 = new_n15857;
  assign po7071 = new_n15858;
  assign po7072 = new_n15859;
  assign po7073 = new_n15860;
  assign po7074 = new_n15861;
  assign po7075 = new_n15862;
  assign po7076 = new_n15863;
  assign po7077 = new_n15864;
  assign po7078 = new_n15865;
  assign po7079 = new_n15866;
  assign po7080 = new_n15867;
  assign po7081 = new_n15868;
  assign po7082 = new_n15869;
  assign po7083 = new_n15870;
  assign po7084 = new_n15871;
  assign po7085 = new_n15872;
  assign po7086 = new_n15873;
  assign po7087 = new_n15874;
  assign po7088 = new_n15875;
  assign po7089 = new_n15876;
  assign po7090 = new_n15877;
  assign po7091 = new_n15878;
  assign po7092 = new_n15879;
  assign po7093 = new_n15880;
  assign po7094 = new_n15881;
  assign po7095 = new_n15882;
  assign po7096 = new_n15883;
  assign po7097 = new_n15884;
  assign po7098 = new_n15885;
  assign po7099 = new_n15886;
  assign po7100 = new_n15887;
  assign po7101 = new_n15888;
  assign po7102 = new_n15890;
  assign po7103 = new_n15891;
  assign po7104 = new_n15892;
  assign po7105 = new_n15893;
  assign po7106 = new_n15894;
  assign po7107 = new_n15895;
  assign po7108 = new_n15896;
  assign po7109 = new_n15897;
  assign po7110 = new_n15898;
  assign po7111 = new_n15899;
  assign po7112 = new_n15900;
  assign po7113 = new_n15901;
  assign po7114 = new_n15902;
  assign po7115 = new_n15903;
  assign po7116 = new_n15904;
  assign po7117 = new_n15905;
  assign po7118 = new_n15906;
  assign po7119 = new_n15907;
  assign po7120 = new_n15908;
  assign po7121 = new_n15909;
  assign po7122 = new_n15910;
  assign po7123 = new_n15911;
  assign po7124 = new_n15912;
  assign po7125 = new_n15913;
  assign po7126 = new_n15914;
  assign po7127 = new_n15915;
  assign po7128 = new_n15916;
  assign po7129 = new_n15917;
  assign po7130 = new_n15918;
  assign po7131 = new_n15919;
  assign po7132 = new_n15920;
  assign po7133 = new_n15921;
  assign po7134 = new_n15923;
  assign po7135 = new_n15924;
  assign po7136 = new_n15925;
  assign po7137 = new_n15926;
  assign po7138 = new_n15927;
  assign po7139 = new_n15928;
  assign po7140 = new_n15929;
  assign po7141 = new_n15930;
  assign po7142 = new_n15931;
  assign po7143 = new_n15932;
  assign po7144 = new_n15933;
  assign po7145 = new_n15934;
  assign po7146 = new_n15935;
  assign po7147 = new_n15936;
  assign po7148 = new_n15937;
  assign po7149 = new_n15938;
  assign po7150 = new_n15939;
  assign po7151 = new_n15940;
  assign po7152 = new_n15941;
  assign po7153 = new_n15942;
  assign po7154 = new_n15943;
  assign po7155 = new_n15944;
  assign po7156 = new_n15945;
  assign po7157 = new_n15946;
  assign po7158 = new_n15947;
  assign po7159 = new_n15948;
  assign po7160 = new_n15949;
  assign po7161 = new_n15950;
  assign po7162 = new_n15951;
  assign po7163 = new_n15952;
  assign po7164 = new_n15953;
  assign po7165 = new_n15954;
endmodule


