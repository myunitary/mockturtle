module adder_opt(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933;
  assign n257 = x128 ^ x0;
  assign n259 = x0 & x128;
  assign n258 = x129 ^ x1;
  assign n260 = n259 ^ n258;
  assign n264 = x130 ^ x2;
  assign n261 = n259 ^ x129;
  assign n262 = n258 & ~n261;
  assign n263 = n262 ^ x1;
  assign n265 = n264 ^ n263;
  assign n269 = x131 ^ x3;
  assign n266 = n263 ^ x130;
  assign n267 = n264 & ~n266;
  assign n268 = n267 ^ x2;
  assign n270 = n269 ^ n268;
  assign n274 = x132 ^ x4;
  assign n271 = n268 ^ x131;
  assign n272 = n269 & ~n271;
  assign n273 = n272 ^ x3;
  assign n275 = n274 ^ n273;
  assign n280 = x133 ^ x5;
  assign n276 = x132 ^ x3;
  assign n277 = n276 ^ n272;
  assign n278 = n274 & ~n277;
  assign n279 = n278 ^ x4;
  assign n281 = n280 ^ n279;
  assign n285 = x134 ^ x6;
  assign n282 = n279 ^ x133;
  assign n283 = n280 & ~n282;
  assign n284 = n283 ^ x5;
  assign n286 = n285 ^ n284;
  assign n291 = x135 ^ x7;
  assign n287 = x134 ^ x5;
  assign n288 = n287 ^ n283;
  assign n289 = n285 & ~n288;
  assign n290 = n289 ^ x6;
  assign n292 = n291 ^ n290;
  assign n296 = x136 ^ x8;
  assign n293 = n290 ^ x135;
  assign n294 = n291 & ~n293;
  assign n295 = n294 ^ x7;
  assign n297 = n296 ^ n295;
  assign n302 = x137 ^ x9;
  assign n298 = x136 ^ x7;
  assign n299 = n298 ^ n294;
  assign n300 = n296 & ~n299;
  assign n301 = n300 ^ x8;
  assign n303 = n302 ^ n301;
  assign n305 = n301 ^ x137;
  assign n306 = n302 & ~n305;
  assign n307 = n306 ^ x9;
  assign n304 = x138 ^ x10;
  assign n308 = n307 ^ n304;
  assign n312 = x139 ^ x11;
  assign n309 = n307 ^ x138;
  assign n310 = n304 & ~n309;
  assign n311 = n310 ^ x10;
  assign n313 = n312 ^ n311;
  assign n317 = x140 ^ x12;
  assign n314 = n311 ^ x139;
  assign n315 = n312 & ~n314;
  assign n316 = n315 ^ x11;
  assign n318 = n317 ^ n316;
  assign n323 = x141 ^ x13;
  assign n319 = x140 ^ x11;
  assign n320 = n319 ^ n315;
  assign n321 = n317 & ~n320;
  assign n322 = n321 ^ x12;
  assign n324 = n323 ^ n322;
  assign n328 = x142 ^ x14;
  assign n325 = n322 ^ x141;
  assign n326 = n323 & ~n325;
  assign n327 = n326 ^ x13;
  assign n329 = n328 ^ n327;
  assign n334 = x143 ^ x15;
  assign n330 = x142 ^ x13;
  assign n331 = n330 ^ n326;
  assign n332 = n328 & ~n331;
  assign n333 = n332 ^ x14;
  assign n335 = n334 ^ n333;
  assign n339 = x144 ^ x16;
  assign n336 = n333 ^ x143;
  assign n337 = n334 & ~n336;
  assign n338 = n337 ^ x15;
  assign n340 = n339 ^ n338;
  assign n345 = x145 ^ x17;
  assign n341 = x144 ^ x15;
  assign n342 = n341 ^ n337;
  assign n343 = n339 & ~n342;
  assign n344 = n343 ^ x16;
  assign n346 = n345 ^ n344;
  assign n350 = x146 ^ x18;
  assign n347 = n344 ^ x145;
  assign n348 = n345 & ~n347;
  assign n349 = n348 ^ x17;
  assign n351 = n350 ^ n349;
  assign n356 = x147 ^ x19;
  assign n352 = x146 ^ x17;
  assign n353 = n352 ^ n348;
  assign n354 = n350 & ~n353;
  assign n355 = n354 ^ x18;
  assign n357 = n356 ^ n355;
  assign n359 = n355 ^ x147;
  assign n360 = n356 & ~n359;
  assign n361 = n360 ^ x19;
  assign n358 = x148 ^ x20;
  assign n362 = n361 ^ n358;
  assign n366 = x149 ^ x21;
  assign n363 = n361 ^ x148;
  assign n364 = n358 & ~n363;
  assign n365 = n364 ^ x20;
  assign n367 = n366 ^ n365;
  assign n371 = x150 ^ x22;
  assign n368 = n365 ^ x149;
  assign n369 = n366 & ~n368;
  assign n370 = n369 ^ x21;
  assign n372 = n371 ^ n370;
  assign n377 = x151 ^ x23;
  assign n373 = x150 ^ x21;
  assign n374 = n373 ^ n369;
  assign n375 = n371 & ~n374;
  assign n376 = n375 ^ x22;
  assign n378 = n377 ^ n376;
  assign n382 = x152 ^ x24;
  assign n379 = n376 ^ x151;
  assign n380 = n377 & ~n379;
  assign n381 = n380 ^ x23;
  assign n383 = n382 ^ n381;
  assign n388 = x153 ^ x25;
  assign n384 = x152 ^ x23;
  assign n385 = n384 ^ n380;
  assign n386 = n382 & ~n385;
  assign n387 = n386 ^ x24;
  assign n389 = n388 ^ n387;
  assign n393 = x154 ^ x26;
  assign n390 = n387 ^ x153;
  assign n391 = n388 & ~n390;
  assign n392 = n391 ^ x25;
  assign n394 = n393 ^ n392;
  assign n399 = x155 ^ x27;
  assign n395 = x154 ^ x25;
  assign n396 = n395 ^ n391;
  assign n397 = n393 & ~n396;
  assign n398 = n397 ^ x26;
  assign n400 = n399 ^ n398;
  assign n404 = x156 ^ x28;
  assign n401 = n398 ^ x155;
  assign n402 = n399 & ~n401;
  assign n403 = n402 ^ x27;
  assign n405 = n404 ^ n403;
  assign n410 = x157 ^ x29;
  assign n406 = x156 ^ x27;
  assign n407 = n406 ^ n402;
  assign n408 = n404 & ~n407;
  assign n409 = n408 ^ x28;
  assign n411 = n410 ^ n409;
  assign n413 = n409 ^ x157;
  assign n414 = n410 & ~n413;
  assign n415 = n414 ^ x29;
  assign n412 = x158 ^ x30;
  assign n416 = n415 ^ n412;
  assign n420 = x159 ^ x31;
  assign n417 = n415 ^ x158;
  assign n418 = n412 & ~n417;
  assign n419 = n418 ^ x30;
  assign n421 = n420 ^ n419;
  assign n425 = x160 ^ x32;
  assign n422 = n419 ^ x159;
  assign n423 = n420 & ~n422;
  assign n424 = n423 ^ x31;
  assign n426 = n425 ^ n424;
  assign n431 = x161 ^ x33;
  assign n427 = x160 ^ x31;
  assign n428 = n427 ^ n423;
  assign n429 = n425 & ~n428;
  assign n430 = n429 ^ x32;
  assign n432 = n431 ^ n430;
  assign n436 = x162 ^ x34;
  assign n433 = n430 ^ x161;
  assign n434 = n431 & ~n433;
  assign n435 = n434 ^ x33;
  assign n437 = n436 ^ n435;
  assign n442 = x163 ^ x35;
  assign n438 = x162 ^ x33;
  assign n439 = n438 ^ n434;
  assign n440 = n436 & ~n439;
  assign n441 = n440 ^ x34;
  assign n443 = n442 ^ n441;
  assign n447 = x164 ^ x36;
  assign n444 = n441 ^ x163;
  assign n445 = n442 & ~n444;
  assign n446 = n445 ^ x35;
  assign n448 = n447 ^ n446;
  assign n453 = x165 ^ x37;
  assign n449 = x164 ^ x35;
  assign n450 = n449 ^ n445;
  assign n451 = n447 & ~n450;
  assign n452 = n451 ^ x36;
  assign n454 = n453 ^ n452;
  assign n458 = x166 ^ x38;
  assign n455 = n452 ^ x165;
  assign n456 = n453 & ~n455;
  assign n457 = n456 ^ x37;
  assign n459 = n458 ^ n457;
  assign n464 = x167 ^ x39;
  assign n460 = x166 ^ x37;
  assign n461 = n460 ^ n456;
  assign n462 = n458 & ~n461;
  assign n463 = n462 ^ x38;
  assign n465 = n464 ^ n463;
  assign n467 = n463 ^ x167;
  assign n468 = n464 & ~n467;
  assign n469 = n468 ^ x39;
  assign n466 = x168 ^ x40;
  assign n470 = n469 ^ n466;
  assign n474 = x169 ^ x41;
  assign n471 = n469 ^ x168;
  assign n472 = n466 & ~n471;
  assign n473 = n472 ^ x40;
  assign n475 = n474 ^ n473;
  assign n479 = x170 ^ x42;
  assign n476 = n473 ^ x169;
  assign n477 = n474 & ~n476;
  assign n478 = n477 ^ x41;
  assign n480 = n479 ^ n478;
  assign n485 = x171 ^ x43;
  assign n481 = x170 ^ x41;
  assign n482 = n481 ^ n477;
  assign n483 = n479 & ~n482;
  assign n484 = n483 ^ x42;
  assign n486 = n485 ^ n484;
  assign n490 = x172 ^ x44;
  assign n487 = n484 ^ x171;
  assign n488 = n485 & ~n487;
  assign n489 = n488 ^ x43;
  assign n491 = n490 ^ n489;
  assign n496 = x173 ^ x45;
  assign n492 = x172 ^ x43;
  assign n493 = n492 ^ n488;
  assign n494 = n490 & ~n493;
  assign n495 = n494 ^ x44;
  assign n497 = n496 ^ n495;
  assign n501 = x174 ^ x46;
  assign n498 = n495 ^ x173;
  assign n499 = n496 & ~n498;
  assign n500 = n499 ^ x45;
  assign n502 = n501 ^ n500;
  assign n507 = x175 ^ x47;
  assign n503 = x174 ^ x45;
  assign n504 = n503 ^ n499;
  assign n505 = n501 & ~n504;
  assign n506 = n505 ^ x46;
  assign n508 = n507 ^ n506;
  assign n512 = x176 ^ x48;
  assign n509 = n506 ^ x175;
  assign n510 = n507 & ~n509;
  assign n511 = n510 ^ x47;
  assign n513 = n512 ^ n511;
  assign n518 = x177 ^ x49;
  assign n514 = x176 ^ x47;
  assign n515 = n514 ^ n510;
  assign n516 = n512 & ~n515;
  assign n517 = n516 ^ x48;
  assign n519 = n518 ^ n517;
  assign n521 = n517 ^ x177;
  assign n522 = n518 & ~n521;
  assign n523 = n522 ^ x49;
  assign n520 = x178 ^ x50;
  assign n524 = n523 ^ n520;
  assign n528 = x179 ^ x51;
  assign n525 = n523 ^ x178;
  assign n526 = n520 & ~n525;
  assign n527 = n526 ^ x50;
  assign n529 = n528 ^ n527;
  assign n533 = x180 ^ x52;
  assign n530 = n527 ^ x179;
  assign n531 = n528 & ~n530;
  assign n532 = n531 ^ x51;
  assign n534 = n533 ^ n532;
  assign n539 = x181 ^ x53;
  assign n535 = x180 ^ x51;
  assign n536 = n535 ^ n531;
  assign n537 = n533 & ~n536;
  assign n538 = n537 ^ x52;
  assign n540 = n539 ^ n538;
  assign n544 = x182 ^ x54;
  assign n541 = n538 ^ x181;
  assign n542 = n539 & ~n541;
  assign n543 = n542 ^ x53;
  assign n545 = n544 ^ n543;
  assign n550 = x183 ^ x55;
  assign n546 = x182 ^ x53;
  assign n547 = n546 ^ n542;
  assign n548 = n544 & ~n547;
  assign n549 = n548 ^ x54;
  assign n551 = n550 ^ n549;
  assign n555 = x184 ^ x56;
  assign n552 = n549 ^ x183;
  assign n553 = n550 & ~n552;
  assign n554 = n553 ^ x55;
  assign n556 = n555 ^ n554;
  assign n561 = x185 ^ x57;
  assign n557 = x184 ^ x55;
  assign n558 = n557 ^ n553;
  assign n559 = n555 & ~n558;
  assign n560 = n559 ^ x56;
  assign n562 = n561 ^ n560;
  assign n566 = x186 ^ x58;
  assign n563 = n560 ^ x185;
  assign n564 = n561 & ~n563;
  assign n565 = n564 ^ x57;
  assign n567 = n566 ^ n565;
  assign n572 = x187 ^ x59;
  assign n568 = x186 ^ x57;
  assign n569 = n568 ^ n564;
  assign n570 = n566 & ~n569;
  assign n571 = n570 ^ x58;
  assign n573 = n572 ^ n571;
  assign n575 = n571 ^ x187;
  assign n576 = n572 & ~n575;
  assign n577 = n576 ^ x59;
  assign n574 = x188 ^ x60;
  assign n578 = n577 ^ n574;
  assign n582 = x189 ^ x61;
  assign n579 = n577 ^ x188;
  assign n580 = n574 & ~n579;
  assign n581 = n580 ^ x60;
  assign n583 = n582 ^ n581;
  assign n587 = x190 ^ x62;
  assign n584 = n581 ^ x189;
  assign n585 = n582 & ~n584;
  assign n586 = n585 ^ x61;
  assign n588 = n587 ^ n586;
  assign n593 = x191 ^ x63;
  assign n589 = x190 ^ x61;
  assign n590 = n589 ^ n585;
  assign n591 = n587 & ~n590;
  assign n592 = n591 ^ x62;
  assign n594 = n593 ^ n592;
  assign n598 = x192 ^ x64;
  assign n595 = n592 ^ x191;
  assign n596 = n593 & ~n595;
  assign n597 = n596 ^ x63;
  assign n599 = n598 ^ n597;
  assign n604 = x193 ^ x65;
  assign n600 = x192 ^ x63;
  assign n601 = n600 ^ n596;
  assign n602 = n598 & ~n601;
  assign n603 = n602 ^ x64;
  assign n605 = n604 ^ n603;
  assign n609 = x194 ^ x66;
  assign n606 = n603 ^ x193;
  assign n607 = n604 & ~n606;
  assign n608 = n607 ^ x65;
  assign n610 = n609 ^ n608;
  assign n615 = x195 ^ x67;
  assign n611 = x194 ^ x65;
  assign n612 = n611 ^ n607;
  assign n613 = n609 & ~n612;
  assign n614 = n613 ^ x66;
  assign n616 = n615 ^ n614;
  assign n620 = x196 ^ x68;
  assign n617 = n614 ^ x195;
  assign n618 = n615 & ~n617;
  assign n619 = n618 ^ x67;
  assign n621 = n620 ^ n619;
  assign n626 = x197 ^ x69;
  assign n622 = x196 ^ x67;
  assign n623 = n622 ^ n618;
  assign n624 = n620 & ~n623;
  assign n625 = n624 ^ x68;
  assign n627 = n626 ^ n625;
  assign n629 = n625 ^ x197;
  assign n630 = n626 & ~n629;
  assign n631 = n630 ^ x69;
  assign n628 = x198 ^ x70;
  assign n632 = n631 ^ n628;
  assign n636 = x199 ^ x71;
  assign n633 = n631 ^ x198;
  assign n634 = n628 & ~n633;
  assign n635 = n634 ^ x70;
  assign n637 = n636 ^ n635;
  assign n641 = x200 ^ x72;
  assign n638 = n635 ^ x199;
  assign n639 = n636 & ~n638;
  assign n640 = n639 ^ x71;
  assign n642 = n641 ^ n640;
  assign n647 = x201 ^ x73;
  assign n643 = x200 ^ x71;
  assign n644 = n643 ^ n639;
  assign n645 = n641 & ~n644;
  assign n646 = n645 ^ x72;
  assign n648 = n647 ^ n646;
  assign n652 = x202 ^ x74;
  assign n649 = n646 ^ x201;
  assign n650 = n647 & ~n649;
  assign n651 = n650 ^ x73;
  assign n653 = n652 ^ n651;
  assign n658 = x203 ^ x75;
  assign n654 = x202 ^ x73;
  assign n655 = n654 ^ n650;
  assign n656 = n652 & ~n655;
  assign n657 = n656 ^ x74;
  assign n659 = n658 ^ n657;
  assign n663 = x204 ^ x76;
  assign n660 = n657 ^ x203;
  assign n661 = n658 & ~n660;
  assign n662 = n661 ^ x75;
  assign n664 = n663 ^ n662;
  assign n669 = x205 ^ x77;
  assign n665 = x204 ^ x75;
  assign n666 = n665 ^ n661;
  assign n667 = n663 & ~n666;
  assign n668 = n667 ^ x76;
  assign n670 = n669 ^ n668;
  assign n674 = x206 ^ x78;
  assign n671 = n668 ^ x205;
  assign n672 = n669 & ~n671;
  assign n673 = n672 ^ x77;
  assign n675 = n674 ^ n673;
  assign n680 = x207 ^ x79;
  assign n676 = x206 ^ x77;
  assign n677 = n676 ^ n672;
  assign n678 = n674 & ~n677;
  assign n679 = n678 ^ x78;
  assign n681 = n680 ^ n679;
  assign n683 = n679 ^ x207;
  assign n684 = n680 & ~n683;
  assign n685 = n684 ^ x79;
  assign n682 = x208 ^ x80;
  assign n686 = n685 ^ n682;
  assign n690 = x209 ^ x81;
  assign n687 = n685 ^ x208;
  assign n688 = n682 & ~n687;
  assign n689 = n688 ^ x80;
  assign n691 = n690 ^ n689;
  assign n695 = x210 ^ x82;
  assign n692 = n689 ^ x209;
  assign n693 = n690 & ~n692;
  assign n694 = n693 ^ x81;
  assign n696 = n695 ^ n694;
  assign n701 = x211 ^ x83;
  assign n697 = x210 ^ x81;
  assign n698 = n697 ^ n693;
  assign n699 = n695 & ~n698;
  assign n700 = n699 ^ x82;
  assign n702 = n701 ^ n700;
  assign n706 = x212 ^ x84;
  assign n703 = n700 ^ x211;
  assign n704 = n701 & ~n703;
  assign n705 = n704 ^ x83;
  assign n707 = n706 ^ n705;
  assign n712 = x213 ^ x85;
  assign n708 = x212 ^ x83;
  assign n709 = n708 ^ n704;
  assign n710 = n706 & ~n709;
  assign n711 = n710 ^ x84;
  assign n713 = n712 ^ n711;
  assign n717 = x214 ^ x86;
  assign n714 = n711 ^ x213;
  assign n715 = n712 & ~n714;
  assign n716 = n715 ^ x85;
  assign n718 = n717 ^ n716;
  assign n723 = x215 ^ x87;
  assign n719 = x214 ^ x85;
  assign n720 = n719 ^ n715;
  assign n721 = n717 & ~n720;
  assign n722 = n721 ^ x86;
  assign n724 = n723 ^ n722;
  assign n728 = x216 ^ x88;
  assign n725 = n722 ^ x215;
  assign n726 = n723 & ~n725;
  assign n727 = n726 ^ x87;
  assign n729 = n728 ^ n727;
  assign n734 = x217 ^ x89;
  assign n730 = x216 ^ x87;
  assign n731 = n730 ^ n726;
  assign n732 = n728 & ~n731;
  assign n733 = n732 ^ x88;
  assign n735 = n734 ^ n733;
  assign n737 = n733 ^ x217;
  assign n738 = n734 & ~n737;
  assign n739 = n738 ^ x89;
  assign n736 = x218 ^ x90;
  assign n740 = n739 ^ n736;
  assign n744 = x219 ^ x91;
  assign n741 = n739 ^ x218;
  assign n742 = n736 & ~n741;
  assign n743 = n742 ^ x90;
  assign n745 = n744 ^ n743;
  assign n747 = n743 ^ x219;
  assign n748 = n744 & ~n747;
  assign n749 = n748 ^ x91;
  assign n746 = x220 ^ x92;
  assign n750 = n749 ^ n746;
  assign n754 = x221 ^ x93;
  assign n751 = n749 ^ x220;
  assign n752 = n746 & ~n751;
  assign n753 = n752 ^ x92;
  assign n755 = n754 ^ n753;
  assign n759 = x222 ^ x94;
  assign n756 = n753 ^ x221;
  assign n757 = n754 & ~n756;
  assign n758 = n757 ^ x93;
  assign n760 = n759 ^ n758;
  assign n764 = x223 ^ x95;
  assign n761 = n758 ^ x222;
  assign n762 = n759 & ~n761;
  assign n763 = n762 ^ x94;
  assign n765 = n764 ^ n763;
  assign n769 = x224 ^ x96;
  assign n766 = n763 ^ x223;
  assign n767 = n764 & ~n766;
  assign n768 = n767 ^ x95;
  assign n770 = n769 ^ n768;
  assign n774 = x225 ^ x97;
  assign n771 = n768 ^ x224;
  assign n772 = n769 & ~n771;
  assign n773 = n772 ^ x96;
  assign n775 = n774 ^ n773;
  assign n779 = x226 ^ x98;
  assign n776 = n773 ^ x225;
  assign n777 = n774 & ~n776;
  assign n778 = n777 ^ x97;
  assign n780 = n779 ^ n778;
  assign n785 = x227 ^ x99;
  assign n781 = x226 ^ x97;
  assign n782 = n781 ^ n777;
  assign n783 = n779 & ~n782;
  assign n784 = n783 ^ x98;
  assign n786 = n785 ^ n784;
  assign n790 = x228 ^ x100;
  assign n787 = n784 ^ x227;
  assign n788 = n785 & ~n787;
  assign n789 = n788 ^ x99;
  assign n791 = n790 ^ n789;
  assign n796 = x229 ^ x101;
  assign n792 = x228 ^ x99;
  assign n793 = n792 ^ n788;
  assign n794 = n790 & ~n793;
  assign n795 = n794 ^ x100;
  assign n797 = n796 ^ n795;
  assign n801 = x230 ^ x102;
  assign n798 = n795 ^ x229;
  assign n799 = n796 & ~n798;
  assign n800 = n799 ^ x101;
  assign n802 = n801 ^ n800;
  assign n807 = x231 ^ x103;
  assign n803 = x230 ^ x101;
  assign n804 = n803 ^ n799;
  assign n805 = n801 & ~n804;
  assign n806 = n805 ^ x102;
  assign n808 = n807 ^ n806;
  assign n812 = x232 ^ x104;
  assign n809 = n806 ^ x231;
  assign n810 = n807 & ~n809;
  assign n811 = n810 ^ x103;
  assign n813 = n812 ^ n811;
  assign n817 = x233 ^ x105;
  assign n814 = n811 ^ x232;
  assign n815 = n812 & ~n814;
  assign n816 = n815 ^ x104;
  assign n818 = n817 ^ n816;
  assign n822 = x234 ^ x106;
  assign n819 = n816 ^ x233;
  assign n820 = n817 & ~n819;
  assign n821 = n820 ^ x105;
  assign n823 = n822 ^ n821;
  assign n828 = x235 ^ x107;
  assign n824 = x234 ^ x105;
  assign n825 = n824 ^ n820;
  assign n826 = n822 & ~n825;
  assign n827 = n826 ^ x106;
  assign n829 = n828 ^ n827;
  assign n833 = x236 ^ x108;
  assign n830 = n827 ^ x235;
  assign n831 = n828 & ~n830;
  assign n832 = n831 ^ x107;
  assign n834 = n833 ^ n832;
  assign n838 = x237 ^ x109;
  assign n835 = n832 ^ x236;
  assign n836 = n833 & ~n835;
  assign n837 = n836 ^ x108;
  assign n839 = n838 ^ n837;
  assign n843 = x238 ^ x110;
  assign n840 = n837 ^ x237;
  assign n841 = n838 & ~n840;
  assign n842 = n841 ^ x109;
  assign n844 = n843 ^ n842;
  assign n849 = x239 ^ x111;
  assign n845 = x238 ^ x109;
  assign n846 = n845 ^ n841;
  assign n847 = n843 & ~n846;
  assign n848 = n847 ^ x110;
  assign n850 = n849 ^ n848;
  assign n854 = x240 ^ x112;
  assign n851 = n848 ^ x239;
  assign n852 = n849 & ~n851;
  assign n853 = n852 ^ x111;
  assign n855 = n854 ^ n853;
  assign n859 = x241 ^ x113;
  assign n856 = n853 ^ x240;
  assign n857 = n854 & ~n856;
  assign n858 = n857 ^ x112;
  assign n860 = n859 ^ n858;
  assign n864 = x242 ^ x114;
  assign n861 = n858 ^ x241;
  assign n862 = n859 & ~n861;
  assign n863 = n862 ^ x113;
  assign n865 = n864 ^ n863;
  assign n869 = x243 ^ x115;
  assign n866 = n863 ^ x242;
  assign n867 = n864 & ~n866;
  assign n868 = n867 ^ x114;
  assign n870 = n869 ^ n868;
  assign n874 = x244 ^ x116;
  assign n871 = n868 ^ x243;
  assign n872 = n869 & ~n871;
  assign n873 = n872 ^ x115;
  assign n875 = n874 ^ n873;
  assign n879 = x245 ^ x117;
  assign n876 = n873 ^ x244;
  assign n877 = n874 & ~n876;
  assign n878 = n877 ^ x116;
  assign n880 = n879 ^ n878;
  assign n884 = x246 ^ x118;
  assign n881 = n878 ^ x245;
  assign n882 = n879 & ~n881;
  assign n883 = n882 ^ x117;
  assign n885 = n884 ^ n883;
  assign n889 = x247 ^ x119;
  assign n886 = n883 ^ x246;
  assign n887 = n884 & ~n886;
  assign n888 = n887 ^ x118;
  assign n890 = n889 ^ n888;
  assign n894 = x248 ^ x120;
  assign n891 = n888 ^ x247;
  assign n892 = n889 & ~n891;
  assign n893 = n892 ^ x119;
  assign n895 = n894 ^ n893;
  assign n899 = x249 ^ x121;
  assign n896 = n893 ^ x248;
  assign n897 = n894 & ~n896;
  assign n898 = n897 ^ x120;
  assign n900 = n899 ^ n898;
  assign n904 = x250 ^ x122;
  assign n901 = n898 ^ x249;
  assign n902 = n899 & ~n901;
  assign n903 = n902 ^ x121;
  assign n905 = n904 ^ n903;
  assign n909 = x251 ^ x123;
  assign n906 = n903 ^ x250;
  assign n907 = n904 & ~n906;
  assign n908 = n907 ^ x122;
  assign n910 = n909 ^ n908;
  assign n914 = x252 ^ x124;
  assign n911 = n908 ^ x251;
  assign n912 = n909 & ~n911;
  assign n913 = n912 ^ x123;
  assign n915 = n914 ^ n913;
  assign n919 = x253 ^ x125;
  assign n916 = n913 ^ x252;
  assign n917 = n914 & ~n916;
  assign n918 = n917 ^ x124;
  assign n920 = n919 ^ n918;
  assign n924 = x254 ^ x126;
  assign n921 = n918 ^ x253;
  assign n922 = n919 & ~n921;
  assign n923 = n922 ^ x125;
  assign n925 = n924 ^ n923;
  assign n929 = x255 ^ x127;
  assign n926 = n923 ^ x254;
  assign n927 = n924 & ~n926;
  assign n928 = n927 ^ x126;
  assign n930 = n929 ^ n928;
  assign n931 = n928 ^ x255;
  assign n932 = n929 & ~n931;
  assign n933 = n932 ^ x127;
  assign y0 = n257;
  assign y1 = n260;
  assign y2 = n265;
  assign y3 = n270;
  assign y4 = n275;
  assign y5 = n281;
  assign y6 = n286;
  assign y7 = n292;
  assign y8 = n297;
  assign y9 = n303;
  assign y10 = n308;
  assign y11 = n313;
  assign y12 = n318;
  assign y13 = n324;
  assign y14 = n329;
  assign y15 = n335;
  assign y16 = n340;
  assign y17 = n346;
  assign y18 = n351;
  assign y19 = n357;
  assign y20 = n362;
  assign y21 = n367;
  assign y22 = n372;
  assign y23 = n378;
  assign y24 = n383;
  assign y25 = n389;
  assign y26 = n394;
  assign y27 = n400;
  assign y28 = n405;
  assign y29 = n411;
  assign y30 = n416;
  assign y31 = n421;
  assign y32 = n426;
  assign y33 = n432;
  assign y34 = n437;
  assign y35 = n443;
  assign y36 = n448;
  assign y37 = n454;
  assign y38 = n459;
  assign y39 = n465;
  assign y40 = n470;
  assign y41 = n475;
  assign y42 = n480;
  assign y43 = n486;
  assign y44 = n491;
  assign y45 = n497;
  assign y46 = n502;
  assign y47 = n508;
  assign y48 = n513;
  assign y49 = n519;
  assign y50 = n524;
  assign y51 = n529;
  assign y52 = n534;
  assign y53 = n540;
  assign y54 = n545;
  assign y55 = n551;
  assign y56 = n556;
  assign y57 = n562;
  assign y58 = n567;
  assign y59 = n573;
  assign y60 = n578;
  assign y61 = n583;
  assign y62 = n588;
  assign y63 = n594;
  assign y64 = n599;
  assign y65 = n605;
  assign y66 = n610;
  assign y67 = n616;
  assign y68 = n621;
  assign y69 = n627;
  assign y70 = n632;
  assign y71 = n637;
  assign y72 = n642;
  assign y73 = n648;
  assign y74 = n653;
  assign y75 = n659;
  assign y76 = n664;
  assign y77 = n670;
  assign y78 = n675;
  assign y79 = n681;
  assign y80 = n686;
  assign y81 = n691;
  assign y82 = n696;
  assign y83 = n702;
  assign y84 = n707;
  assign y85 = n713;
  assign y86 = n718;
  assign y87 = n724;
  assign y88 = n729;
  assign y89 = n735;
  assign y90 = n740;
  assign y91 = n745;
  assign y92 = n750;
  assign y93 = n755;
  assign y94 = n760;
  assign y95 = n765;
  assign y96 = n770;
  assign y97 = n775;
  assign y98 = n780;
  assign y99 = n786;
  assign y100 = n791;
  assign y101 = n797;
  assign y102 = n802;
  assign y103 = n808;
  assign y104 = n813;
  assign y105 = n818;
  assign y106 = n823;
  assign y107 = n829;
  assign y108 = n834;
  assign y109 = n839;
  assign y110 = n844;
  assign y111 = n850;
  assign y112 = n855;
  assign y113 = n860;
  assign y114 = n865;
  assign y115 = n870;
  assign y116 = n875;
  assign y117 = n880;
  assign y118 = n885;
  assign y119 = n890;
  assign y120 = n895;
  assign y121 = n900;
  assign y122 = n905;
  assign y123 = n910;
  assign y124 = n915;
  assign y125 = n920;
  assign y126 = n925;
  assign y127 = n930;
  assign y128 = n933;
endmodule
