module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 ;
  assign n84 = x0 & ~x8 ;
  assign n49 = x8 ^ x0 ;
  assign n82 = x1 & ~x9 ;
  assign n83 = ~n49 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n50 = x9 ^ x1 ;
  assign n51 = ~n49 & ~n50 ;
  assign n79 = x2 & ~x10 ;
  assign n52 = x10 ^ x2 ;
  assign n77 = x3 & ~x11 ;
  assign n78 = ~n52 & n77 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n51 & n80 ;
  assign n86 = n85 ^ n81 ;
  assign n53 = x11 ^ x3 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n51 & n54 ;
  assign n73 = x4 & ~x12 ;
  assign n56 = x12 ^ x4 ;
  assign n71 = x5 & ~x13 ;
  assign n72 = ~n56 & n71 ;
  assign n74 = n73 ^ n72 ;
  assign n57 = x13 ^ x5 ;
  assign n58 = ~n56 & ~n57 ;
  assign n68 = x6 & ~x14 ;
  assign n59 = x14 ^ x6 ;
  assign n64 = x7 & x15 ;
  assign n65 = n64 ^ x7 ;
  assign n66 = n59 & n65 ;
  assign n67 = n66 ^ n65 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n58 & n69 ;
  assign n75 = n74 ^ n70 ;
  assign n76 = n55 & n75 ;
  assign n87 = n86 ^ n76 ;
  assign n60 = x15 ^ x7 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 & n62 ;
  assign n88 = n87 ^ n63 ;
  assign n353 = x0 & ~n88 ;
  assign n352 = x8 & n88 ;
  assign n354 = n353 ^ n352 ;
  assign n90 = x8 & ~n88 ;
  assign n89 = x0 & n88 ;
  assign n91 = n90 ^ n89 ;
  assign n149 = ~x16 & n91 ;
  assign n92 = n91 ^ x16 ;
  assign n94 = x9 & ~n88 ;
  assign n93 = x1 & n88 ;
  assign n95 = n94 ^ n93 ;
  assign n147 = ~x17 & n95 ;
  assign n148 = ~n92 & n147 ;
  assign n150 = n149 ^ n148 ;
  assign n96 = n95 ^ x17 ;
  assign n97 = ~n92 & ~n96 ;
  assign n99 = x10 & ~n88 ;
  assign n98 = x2 & n88 ;
  assign n100 = n99 ^ n98 ;
  assign n144 = ~x18 & n100 ;
  assign n101 = n100 ^ x18 ;
  assign n103 = x11 & ~n88 ;
  assign n102 = x3 & n88 ;
  assign n104 = n103 ^ n102 ;
  assign n142 = ~x19 & n104 ;
  assign n143 = ~n101 & n142 ;
  assign n145 = n144 ^ n143 ;
  assign n146 = n97 & n145 ;
  assign n151 = n150 ^ n146 ;
  assign n105 = n104 ^ x19 ;
  assign n106 = ~n101 & ~n105 ;
  assign n107 = n97 & n106 ;
  assign n109 = x12 & ~n88 ;
  assign n108 = x4 & n88 ;
  assign n110 = n109 ^ n108 ;
  assign n138 = ~x20 & n110 ;
  assign n111 = n110 ^ x20 ;
  assign n113 = x13 & ~n88 ;
  assign n112 = x5 & n88 ;
  assign n114 = n113 ^ n112 ;
  assign n136 = ~x21 & n114 ;
  assign n137 = ~n111 & n136 ;
  assign n139 = n138 ^ n137 ;
  assign n115 = n114 ^ x21 ;
  assign n116 = ~n111 & ~n115 ;
  assign n118 = x14 & ~n88 ;
  assign n117 = x6 & n88 ;
  assign n119 = n118 ^ n117 ;
  assign n133 = ~x22 & n119 ;
  assign n120 = n119 ^ x22 ;
  assign n122 = x15 & n88 ;
  assign n123 = n122 ^ x15 ;
  assign n121 = x7 & n88 ;
  assign n124 = n123 ^ n121 ;
  assign n129 = x23 & n124 ;
  assign n130 = n129 ^ n124 ;
  assign n131 = n120 & n130 ;
  assign n132 = n131 ^ n130 ;
  assign n134 = n133 ^ n132 ;
  assign n135 = n116 & n134 ;
  assign n140 = n139 ^ n135 ;
  assign n141 = n107 & n140 ;
  assign n152 = n151 ^ n141 ;
  assign n125 = n124 ^ x23 ;
  assign n126 = ~n120 & ~n125 ;
  assign n127 = n116 & n126 ;
  assign n128 = n107 & n127 ;
  assign n153 = n152 ^ n128 ;
  assign n356 = n91 & ~n153 ;
  assign n355 = x16 & n153 ;
  assign n357 = n356 ^ n355 ;
  assign n433 = n354 & ~n357 ;
  assign n358 = n357 ^ n354 ;
  assign n360 = n95 & ~n153 ;
  assign n359 = x17 & n153 ;
  assign n361 = n360 ^ n359 ;
  assign n363 = x1 & ~n88 ;
  assign n362 = x9 & n88 ;
  assign n364 = n363 ^ n362 ;
  assign n431 = ~n361 & n364 ;
  assign n432 = ~n358 & n431 ;
  assign n434 = n433 ^ n432 ;
  assign n365 = n364 ^ n361 ;
  assign n366 = ~n358 & ~n365 ;
  assign n368 = x2 & ~n88 ;
  assign n367 = x10 & n88 ;
  assign n369 = n368 ^ n367 ;
  assign n371 = n100 & ~n153 ;
  assign n370 = x18 & n153 ;
  assign n372 = n371 ^ n370 ;
  assign n428 = n369 & ~n372 ;
  assign n373 = n372 ^ n369 ;
  assign n375 = x3 & ~n88 ;
  assign n374 = x11 & n88 ;
  assign n376 = n375 ^ n374 ;
  assign n378 = n104 & ~n153 ;
  assign n377 = x19 & n153 ;
  assign n379 = n378 ^ n377 ;
  assign n426 = n376 & ~n379 ;
  assign n427 = ~n373 & n426 ;
  assign n429 = n428 ^ n427 ;
  assign n430 = n366 & n429 ;
  assign n435 = n434 ^ n430 ;
  assign n380 = n379 ^ n376 ;
  assign n381 = ~n373 & ~n380 ;
  assign n382 = n366 & n381 ;
  assign n384 = x4 & ~n88 ;
  assign n383 = x12 & n88 ;
  assign n385 = n384 ^ n383 ;
  assign n387 = n110 & ~n153 ;
  assign n386 = x20 & n153 ;
  assign n388 = n387 ^ n386 ;
  assign n422 = n385 & ~n388 ;
  assign n389 = n388 ^ n385 ;
  assign n391 = x5 & ~n88 ;
  assign n390 = x13 & n88 ;
  assign n392 = n391 ^ n390 ;
  assign n394 = n114 & ~n153 ;
  assign n393 = x21 & n153 ;
  assign n395 = n394 ^ n393 ;
  assign n420 = n392 & ~n395 ;
  assign n421 = ~n389 & n420 ;
  assign n423 = n422 ^ n421 ;
  assign n396 = n395 ^ n392 ;
  assign n397 = ~n389 & ~n396 ;
  assign n399 = x6 & ~n88 ;
  assign n398 = x14 & n88 ;
  assign n400 = n399 ^ n398 ;
  assign n402 = n119 & ~n153 ;
  assign n401 = x22 & n153 ;
  assign n403 = n402 ^ n401 ;
  assign n417 = n400 & ~n403 ;
  assign n404 = n403 ^ n400 ;
  assign n188 = n124 & n153 ;
  assign n405 = n188 ^ n124 ;
  assign n186 = x23 & n153 ;
  assign n406 = n405 ^ n186 ;
  assign n407 = x7 & ~n88 ;
  assign n408 = n407 ^ n122 ;
  assign n413 = n406 & n408 ;
  assign n414 = n413 ^ n408 ;
  assign n415 = n404 & n414 ;
  assign n416 = n415 ^ n414 ;
  assign n418 = n417 ^ n416 ;
  assign n419 = n397 & n418 ;
  assign n424 = n423 ^ n419 ;
  assign n425 = n382 & n424 ;
  assign n436 = n435 ^ n425 ;
  assign n409 = n408 ^ n406 ;
  assign n410 = ~n404 & ~n409 ;
  assign n411 = n397 & n410 ;
  assign n412 = n382 & n411 ;
  assign n437 = n436 ^ n412 ;
  assign n705 = n354 & ~n437 ;
  assign n704 = n357 & n437 ;
  assign n706 = n705 ^ n704 ;
  assign n439 = n357 & ~n437 ;
  assign n438 = n354 & n437 ;
  assign n440 = n439 ^ n438 ;
  assign n155 = x16 & ~n153 ;
  assign n154 = n91 & n153 ;
  assign n156 = n155 ^ n154 ;
  assign n214 = ~x24 & n156 ;
  assign n157 = n156 ^ x24 ;
  assign n159 = x17 & ~n153 ;
  assign n158 = n95 & n153 ;
  assign n160 = n159 ^ n158 ;
  assign n212 = ~x25 & n160 ;
  assign n213 = ~n157 & n212 ;
  assign n215 = n214 ^ n213 ;
  assign n161 = n160 ^ x25 ;
  assign n162 = ~n157 & ~n161 ;
  assign n164 = x18 & ~n153 ;
  assign n163 = n100 & n153 ;
  assign n165 = n164 ^ n163 ;
  assign n209 = ~x26 & n165 ;
  assign n166 = n165 ^ x26 ;
  assign n168 = x19 & ~n153 ;
  assign n167 = n104 & n153 ;
  assign n169 = n168 ^ n167 ;
  assign n207 = ~x27 & n169 ;
  assign n208 = ~n166 & n207 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n162 & n210 ;
  assign n216 = n215 ^ n211 ;
  assign n170 = n169 ^ x27 ;
  assign n171 = ~n166 & ~n170 ;
  assign n172 = n162 & n171 ;
  assign n174 = x20 & ~n153 ;
  assign n173 = n110 & n153 ;
  assign n175 = n174 ^ n173 ;
  assign n203 = ~x28 & n175 ;
  assign n176 = n175 ^ x28 ;
  assign n178 = x21 & ~n153 ;
  assign n177 = n114 & n153 ;
  assign n179 = n178 ^ n177 ;
  assign n201 = ~x29 & n179 ;
  assign n202 = ~n176 & n201 ;
  assign n204 = n203 ^ n202 ;
  assign n180 = n179 ^ x29 ;
  assign n181 = ~n176 & ~n180 ;
  assign n183 = x22 & ~n153 ;
  assign n182 = n119 & n153 ;
  assign n184 = n183 ^ n182 ;
  assign n198 = ~x30 & n184 ;
  assign n185 = n184 ^ x30 ;
  assign n187 = n186 ^ x23 ;
  assign n189 = n188 ^ n187 ;
  assign n194 = x31 & n189 ;
  assign n195 = n194 ^ n189 ;
  assign n196 = n185 & n195 ;
  assign n197 = n196 ^ n195 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = n181 & n199 ;
  assign n205 = n204 ^ n200 ;
  assign n206 = n172 & n205 ;
  assign n217 = n216 ^ n206 ;
  assign n190 = n189 ^ x31 ;
  assign n191 = ~n185 & ~n190 ;
  assign n192 = n181 & n191 ;
  assign n193 = n172 & n192 ;
  assign n218 = n217 ^ n193 ;
  assign n442 = n156 & ~n218 ;
  assign n441 = x24 & n218 ;
  assign n443 = n442 ^ n441 ;
  assign n521 = n440 & ~n443 ;
  assign n444 = n443 ^ n440 ;
  assign n446 = n160 & ~n218 ;
  assign n445 = x25 & n218 ;
  assign n447 = n446 ^ n445 ;
  assign n449 = n361 & ~n437 ;
  assign n448 = n364 & n437 ;
  assign n450 = n449 ^ n448 ;
  assign n519 = ~n447 & n450 ;
  assign n520 = ~n444 & n519 ;
  assign n522 = n521 ^ n520 ;
  assign n451 = n450 ^ n447 ;
  assign n452 = ~n444 & ~n451 ;
  assign n454 = n372 & ~n437 ;
  assign n453 = n369 & n437 ;
  assign n455 = n454 ^ n453 ;
  assign n457 = n165 & ~n218 ;
  assign n456 = x26 & n218 ;
  assign n458 = n457 ^ n456 ;
  assign n516 = n455 & ~n458 ;
  assign n459 = n458 ^ n455 ;
  assign n461 = n379 & ~n437 ;
  assign n460 = n376 & n437 ;
  assign n462 = n461 ^ n460 ;
  assign n464 = n169 & ~n218 ;
  assign n463 = x27 & n218 ;
  assign n465 = n464 ^ n463 ;
  assign n514 = n462 & ~n465 ;
  assign n515 = ~n459 & n514 ;
  assign n517 = n516 ^ n515 ;
  assign n518 = n452 & n517 ;
  assign n523 = n522 ^ n518 ;
  assign n466 = n465 ^ n462 ;
  assign n467 = ~n459 & ~n466 ;
  assign n468 = n452 & n467 ;
  assign n470 = n388 & ~n437 ;
  assign n469 = n385 & n437 ;
  assign n471 = n470 ^ n469 ;
  assign n473 = n175 & ~n218 ;
  assign n472 = x28 & n218 ;
  assign n474 = n473 ^ n472 ;
  assign n510 = n471 & ~n474 ;
  assign n475 = n474 ^ n471 ;
  assign n477 = n395 & ~n437 ;
  assign n476 = n392 & n437 ;
  assign n478 = n477 ^ n476 ;
  assign n480 = n179 & ~n218 ;
  assign n479 = x29 & n218 ;
  assign n481 = n480 ^ n479 ;
  assign n508 = n478 & ~n481 ;
  assign n509 = ~n475 & n508 ;
  assign n511 = n510 ^ n509 ;
  assign n482 = n481 ^ n478 ;
  assign n483 = ~n475 & ~n482 ;
  assign n485 = n403 & ~n437 ;
  assign n484 = n400 & n437 ;
  assign n486 = n485 ^ n484 ;
  assign n488 = n184 & ~n218 ;
  assign n487 = x30 & n218 ;
  assign n489 = n488 ^ n487 ;
  assign n505 = n486 & ~n489 ;
  assign n490 = n489 ^ n486 ;
  assign n253 = n189 & n218 ;
  assign n491 = n253 ^ n189 ;
  assign n251 = x31 & n218 ;
  assign n492 = n491 ^ n251 ;
  assign n494 = n406 & n437 ;
  assign n495 = n494 ^ n406 ;
  assign n493 = n408 & n437 ;
  assign n496 = n495 ^ n493 ;
  assign n501 = n492 & n496 ;
  assign n502 = n501 ^ n496 ;
  assign n503 = n490 & n502 ;
  assign n504 = n503 ^ n502 ;
  assign n506 = n505 ^ n504 ;
  assign n507 = n483 & n506 ;
  assign n512 = n511 ^ n507 ;
  assign n513 = n468 & n512 ;
  assign n524 = n523 ^ n513 ;
  assign n497 = n496 ^ n492 ;
  assign n498 = ~n490 & ~n497 ;
  assign n499 = n483 & n498 ;
  assign n500 = n468 & n499 ;
  assign n525 = n524 ^ n500 ;
  assign n708 = n440 & ~n525 ;
  assign n707 = n443 & n525 ;
  assign n709 = n708 ^ n707 ;
  assign n785 = n706 & ~n709 ;
  assign n710 = n709 ^ n706 ;
  assign n712 = n450 & ~n525 ;
  assign n711 = n447 & n525 ;
  assign n713 = n712 ^ n711 ;
  assign n715 = n364 & ~n437 ;
  assign n714 = n361 & n437 ;
  assign n716 = n715 ^ n714 ;
  assign n783 = ~n713 & n716 ;
  assign n784 = ~n710 & n783 ;
  assign n786 = n785 ^ n784 ;
  assign n717 = n716 ^ n713 ;
  assign n718 = ~n710 & ~n717 ;
  assign n720 = n369 & ~n437 ;
  assign n719 = n372 & n437 ;
  assign n721 = n720 ^ n719 ;
  assign n723 = n455 & ~n525 ;
  assign n722 = n458 & n525 ;
  assign n724 = n723 ^ n722 ;
  assign n780 = n721 & ~n724 ;
  assign n725 = n724 ^ n721 ;
  assign n727 = n376 & ~n437 ;
  assign n726 = n379 & n437 ;
  assign n728 = n727 ^ n726 ;
  assign n730 = n462 & ~n525 ;
  assign n729 = n465 & n525 ;
  assign n731 = n730 ^ n729 ;
  assign n778 = n728 & ~n731 ;
  assign n779 = ~n725 & n778 ;
  assign n781 = n780 ^ n779 ;
  assign n782 = n718 & n781 ;
  assign n787 = n786 ^ n782 ;
  assign n732 = n731 ^ n728 ;
  assign n733 = ~n725 & ~n732 ;
  assign n734 = n718 & n733 ;
  assign n736 = n385 & ~n437 ;
  assign n735 = n388 & n437 ;
  assign n737 = n736 ^ n735 ;
  assign n739 = n471 & ~n525 ;
  assign n738 = n474 & n525 ;
  assign n740 = n739 ^ n738 ;
  assign n774 = n737 & ~n740 ;
  assign n741 = n740 ^ n737 ;
  assign n743 = n392 & ~n437 ;
  assign n742 = n395 & n437 ;
  assign n744 = n743 ^ n742 ;
  assign n746 = n478 & ~n525 ;
  assign n745 = n481 & n525 ;
  assign n747 = n746 ^ n745 ;
  assign n772 = n744 & ~n747 ;
  assign n773 = ~n741 & n772 ;
  assign n775 = n774 ^ n773 ;
  assign n748 = n747 ^ n744 ;
  assign n749 = ~n741 & ~n748 ;
  assign n751 = n400 & ~n437 ;
  assign n750 = n403 & n437 ;
  assign n752 = n751 ^ n750 ;
  assign n754 = n486 & ~n525 ;
  assign n753 = n489 & n525 ;
  assign n755 = n754 ^ n753 ;
  assign n769 = n752 & ~n755 ;
  assign n756 = n755 ^ n752 ;
  assign n583 = n496 & n525 ;
  assign n757 = n583 ^ n496 ;
  assign n581 = n492 & n525 ;
  assign n758 = n757 ^ n581 ;
  assign n759 = n408 & ~n437 ;
  assign n760 = n759 ^ n494 ;
  assign n765 = n758 & n760 ;
  assign n766 = n765 ^ n760 ;
  assign n767 = n756 & n766 ;
  assign n768 = n767 ^ n766 ;
  assign n770 = n769 ^ n768 ;
  assign n771 = n749 & n770 ;
  assign n776 = n775 ^ n771 ;
  assign n777 = n734 & n776 ;
  assign n788 = n787 ^ n777 ;
  assign n761 = n760 ^ n758 ;
  assign n762 = ~n756 & ~n761 ;
  assign n763 = n749 & n762 ;
  assign n764 = n734 & n763 ;
  assign n789 = n788 ^ n764 ;
  assign n969 = n706 & ~n789 ;
  assign n968 = n709 & n789 ;
  assign n970 = n969 ^ n968 ;
  assign n791 = n709 & ~n789 ;
  assign n790 = n706 & n789 ;
  assign n792 = n791 ^ n790 ;
  assign n527 = n443 & ~n525 ;
  assign n526 = n440 & n525 ;
  assign n528 = n527 ^ n526 ;
  assign n220 = x24 & ~n218 ;
  assign n219 = n156 & n218 ;
  assign n221 = n220 ^ n219 ;
  assign n279 = ~x32 & n221 ;
  assign n222 = n221 ^ x32 ;
  assign n224 = x25 & ~n218 ;
  assign n223 = n160 & n218 ;
  assign n225 = n224 ^ n223 ;
  assign n277 = ~x33 & n225 ;
  assign n278 = ~n222 & n277 ;
  assign n280 = n279 ^ n278 ;
  assign n226 = n225 ^ x33 ;
  assign n227 = ~n222 & ~n226 ;
  assign n229 = x26 & ~n218 ;
  assign n228 = n165 & n218 ;
  assign n230 = n229 ^ n228 ;
  assign n274 = ~x34 & n230 ;
  assign n231 = n230 ^ x34 ;
  assign n233 = x27 & ~n218 ;
  assign n232 = n169 & n218 ;
  assign n234 = n233 ^ n232 ;
  assign n272 = ~x35 & n234 ;
  assign n273 = ~n231 & n272 ;
  assign n275 = n274 ^ n273 ;
  assign n276 = n227 & n275 ;
  assign n281 = n280 ^ n276 ;
  assign n235 = n234 ^ x35 ;
  assign n236 = ~n231 & ~n235 ;
  assign n237 = n227 & n236 ;
  assign n239 = x28 & ~n218 ;
  assign n238 = n175 & n218 ;
  assign n240 = n239 ^ n238 ;
  assign n268 = ~x36 & n240 ;
  assign n241 = n240 ^ x36 ;
  assign n243 = x29 & ~n218 ;
  assign n242 = n179 & n218 ;
  assign n244 = n243 ^ n242 ;
  assign n266 = ~x37 & n244 ;
  assign n267 = ~n241 & n266 ;
  assign n269 = n268 ^ n267 ;
  assign n245 = n244 ^ x37 ;
  assign n246 = ~n241 & ~n245 ;
  assign n248 = x30 & ~n218 ;
  assign n247 = n184 & n218 ;
  assign n249 = n248 ^ n247 ;
  assign n263 = ~x38 & n249 ;
  assign n250 = n249 ^ x38 ;
  assign n252 = n251 ^ x31 ;
  assign n254 = n253 ^ n252 ;
  assign n259 = x39 & n254 ;
  assign n260 = n259 ^ n254 ;
  assign n261 = n250 & n260 ;
  assign n262 = n261 ^ n260 ;
  assign n264 = n263 ^ n262 ;
  assign n265 = n246 & n264 ;
  assign n270 = n269 ^ n265 ;
  assign n271 = n237 & n270 ;
  assign n282 = n281 ^ n271 ;
  assign n255 = n254 ^ x39 ;
  assign n256 = ~n250 & ~n255 ;
  assign n257 = n246 & n256 ;
  assign n258 = n237 & n257 ;
  assign n283 = n282 ^ n258 ;
  assign n530 = n221 & ~n283 ;
  assign n529 = x32 & n283 ;
  assign n531 = n530 ^ n529 ;
  assign n609 = n528 & ~n531 ;
  assign n532 = n531 ^ n528 ;
  assign n534 = n225 & ~n283 ;
  assign n533 = x33 & n283 ;
  assign n535 = n534 ^ n533 ;
  assign n537 = n447 & ~n525 ;
  assign n536 = n450 & n525 ;
  assign n538 = n537 ^ n536 ;
  assign n607 = ~n535 & n538 ;
  assign n608 = ~n532 & n607 ;
  assign n610 = n609 ^ n608 ;
  assign n539 = n538 ^ n535 ;
  assign n540 = ~n532 & ~n539 ;
  assign n542 = n458 & ~n525 ;
  assign n541 = n455 & n525 ;
  assign n543 = n542 ^ n541 ;
  assign n545 = n230 & ~n283 ;
  assign n544 = x34 & n283 ;
  assign n546 = n545 ^ n544 ;
  assign n604 = n543 & ~n546 ;
  assign n547 = n546 ^ n543 ;
  assign n549 = n465 & ~n525 ;
  assign n548 = n462 & n525 ;
  assign n550 = n549 ^ n548 ;
  assign n552 = n234 & ~n283 ;
  assign n551 = x35 & n283 ;
  assign n553 = n552 ^ n551 ;
  assign n602 = n550 & ~n553 ;
  assign n603 = ~n547 & n602 ;
  assign n605 = n604 ^ n603 ;
  assign n606 = n540 & n605 ;
  assign n611 = n610 ^ n606 ;
  assign n554 = n553 ^ n550 ;
  assign n555 = ~n547 & ~n554 ;
  assign n556 = n540 & n555 ;
  assign n558 = n474 & ~n525 ;
  assign n557 = n471 & n525 ;
  assign n559 = n558 ^ n557 ;
  assign n561 = n240 & ~n283 ;
  assign n560 = x36 & n283 ;
  assign n562 = n561 ^ n560 ;
  assign n598 = n559 & ~n562 ;
  assign n563 = n562 ^ n559 ;
  assign n565 = n481 & ~n525 ;
  assign n564 = n478 & n525 ;
  assign n566 = n565 ^ n564 ;
  assign n568 = n244 & ~n283 ;
  assign n567 = x37 & n283 ;
  assign n569 = n568 ^ n567 ;
  assign n596 = n566 & ~n569 ;
  assign n597 = ~n563 & n596 ;
  assign n599 = n598 ^ n597 ;
  assign n570 = n569 ^ n566 ;
  assign n571 = ~n563 & ~n570 ;
  assign n573 = n489 & ~n525 ;
  assign n572 = n486 & n525 ;
  assign n574 = n573 ^ n572 ;
  assign n576 = n249 & ~n283 ;
  assign n575 = x38 & n283 ;
  assign n577 = n576 ^ n575 ;
  assign n593 = n574 & ~n577 ;
  assign n578 = n577 ^ n574 ;
  assign n318 = n254 & n283 ;
  assign n579 = n318 ^ n254 ;
  assign n316 = x39 & n283 ;
  assign n580 = n579 ^ n316 ;
  assign n582 = n581 ^ n492 ;
  assign n584 = n583 ^ n582 ;
  assign n589 = n580 & n584 ;
  assign n590 = n589 ^ n584 ;
  assign n591 = n578 & n590 ;
  assign n592 = n591 ^ n590 ;
  assign n594 = n593 ^ n592 ;
  assign n595 = n571 & n594 ;
  assign n600 = n599 ^ n595 ;
  assign n601 = n556 & n600 ;
  assign n612 = n611 ^ n601 ;
  assign n585 = n584 ^ n580 ;
  assign n586 = ~n578 & ~n585 ;
  assign n587 = n571 & n586 ;
  assign n588 = n556 & n587 ;
  assign n613 = n612 ^ n588 ;
  assign n794 = n528 & ~n613 ;
  assign n793 = n531 & n613 ;
  assign n795 = n794 ^ n793 ;
  assign n873 = n792 & ~n795 ;
  assign n796 = n795 ^ n792 ;
  assign n798 = n538 & ~n613 ;
  assign n797 = n535 & n613 ;
  assign n799 = n798 ^ n797 ;
  assign n801 = n713 & ~n789 ;
  assign n800 = n716 & n789 ;
  assign n802 = n801 ^ n800 ;
  assign n871 = ~n799 & n802 ;
  assign n872 = ~n796 & n871 ;
  assign n874 = n873 ^ n872 ;
  assign n803 = n802 ^ n799 ;
  assign n804 = ~n796 & ~n803 ;
  assign n806 = n724 & ~n789 ;
  assign n805 = n721 & n789 ;
  assign n807 = n806 ^ n805 ;
  assign n809 = n543 & ~n613 ;
  assign n808 = n546 & n613 ;
  assign n810 = n809 ^ n808 ;
  assign n868 = n807 & ~n810 ;
  assign n811 = n810 ^ n807 ;
  assign n813 = n731 & ~n789 ;
  assign n812 = n728 & n789 ;
  assign n814 = n813 ^ n812 ;
  assign n816 = n550 & ~n613 ;
  assign n815 = n553 & n613 ;
  assign n817 = n816 ^ n815 ;
  assign n866 = n814 & ~n817 ;
  assign n867 = ~n811 & n866 ;
  assign n869 = n868 ^ n867 ;
  assign n870 = n804 & n869 ;
  assign n875 = n874 ^ n870 ;
  assign n818 = n817 ^ n814 ;
  assign n819 = ~n811 & ~n818 ;
  assign n820 = n804 & n819 ;
  assign n822 = n740 & ~n789 ;
  assign n821 = n737 & n789 ;
  assign n823 = n822 ^ n821 ;
  assign n825 = n559 & ~n613 ;
  assign n824 = n562 & n613 ;
  assign n826 = n825 ^ n824 ;
  assign n862 = n823 & ~n826 ;
  assign n827 = n826 ^ n823 ;
  assign n829 = n747 & ~n789 ;
  assign n828 = n744 & n789 ;
  assign n830 = n829 ^ n828 ;
  assign n832 = n566 & ~n613 ;
  assign n831 = n569 & n613 ;
  assign n833 = n832 ^ n831 ;
  assign n860 = n830 & ~n833 ;
  assign n861 = ~n827 & n860 ;
  assign n863 = n862 ^ n861 ;
  assign n834 = n833 ^ n830 ;
  assign n835 = ~n827 & ~n834 ;
  assign n837 = n755 & ~n789 ;
  assign n836 = n752 & n789 ;
  assign n838 = n837 ^ n836 ;
  assign n840 = n574 & ~n613 ;
  assign n839 = n577 & n613 ;
  assign n841 = n840 ^ n839 ;
  assign n857 = n838 & ~n841 ;
  assign n842 = n841 ^ n838 ;
  assign n666 = n584 & n613 ;
  assign n843 = n666 ^ n584 ;
  assign n664 = n580 & n613 ;
  assign n844 = n843 ^ n664 ;
  assign n846 = n758 & n789 ;
  assign n847 = n846 ^ n758 ;
  assign n845 = n760 & n789 ;
  assign n848 = n847 ^ n845 ;
  assign n853 = n844 & n848 ;
  assign n854 = n853 ^ n848 ;
  assign n855 = n842 & n854 ;
  assign n856 = n855 ^ n854 ;
  assign n858 = n857 ^ n856 ;
  assign n859 = n835 & n858 ;
  assign n864 = n863 ^ n859 ;
  assign n865 = n820 & n864 ;
  assign n876 = n875 ^ n865 ;
  assign n849 = n848 ^ n844 ;
  assign n850 = ~n842 & ~n849 ;
  assign n851 = n835 & n850 ;
  assign n852 = n820 & n851 ;
  assign n877 = n876 ^ n852 ;
  assign n972 = n792 & ~n877 ;
  assign n971 = n795 & n877 ;
  assign n973 = n972 ^ n971 ;
  assign n1049 = n970 & ~n973 ;
  assign n974 = n973 ^ n970 ;
  assign n976 = n802 & ~n877 ;
  assign n975 = n799 & n877 ;
  assign n977 = n976 ^ n975 ;
  assign n979 = n716 & ~n789 ;
  assign n978 = n713 & n789 ;
  assign n980 = n979 ^ n978 ;
  assign n1047 = ~n977 & n980 ;
  assign n1048 = ~n974 & n1047 ;
  assign n1050 = n1049 ^ n1048 ;
  assign n981 = n980 ^ n977 ;
  assign n982 = ~n974 & ~n981 ;
  assign n984 = n721 & ~n789 ;
  assign n983 = n724 & n789 ;
  assign n985 = n984 ^ n983 ;
  assign n987 = n807 & ~n877 ;
  assign n986 = n810 & n877 ;
  assign n988 = n987 ^ n986 ;
  assign n1044 = n985 & ~n988 ;
  assign n989 = n988 ^ n985 ;
  assign n991 = n728 & ~n789 ;
  assign n990 = n731 & n789 ;
  assign n992 = n991 ^ n990 ;
  assign n994 = n814 & ~n877 ;
  assign n993 = n817 & n877 ;
  assign n995 = n994 ^ n993 ;
  assign n1042 = n992 & ~n995 ;
  assign n1043 = ~n989 & n1042 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n1046 = n982 & n1045 ;
  assign n1051 = n1050 ^ n1046 ;
  assign n996 = n995 ^ n992 ;
  assign n997 = ~n989 & ~n996 ;
  assign n998 = n982 & n997 ;
  assign n1000 = n737 & ~n789 ;
  assign n999 = n740 & n789 ;
  assign n1001 = n1000 ^ n999 ;
  assign n1003 = n823 & ~n877 ;
  assign n1002 = n826 & n877 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1038 = n1001 & ~n1004 ;
  assign n1005 = n1004 ^ n1001 ;
  assign n1007 = n744 & ~n789 ;
  assign n1006 = n747 & n789 ;
  assign n1008 = n1007 ^ n1006 ;
  assign n1010 = n830 & ~n877 ;
  assign n1009 = n833 & n877 ;
  assign n1011 = n1010 ^ n1009 ;
  assign n1036 = n1008 & ~n1011 ;
  assign n1037 = ~n1005 & n1036 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1012 = n1011 ^ n1008 ;
  assign n1013 = ~n1005 & ~n1012 ;
  assign n1015 = n752 & ~n789 ;
  assign n1014 = n755 & n789 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1018 = n838 & ~n877 ;
  assign n1017 = n841 & n877 ;
  assign n1019 = n1018 ^ n1017 ;
  assign n1033 = n1016 & ~n1019 ;
  assign n1020 = n1019 ^ n1016 ;
  assign n930 = n848 & n877 ;
  assign n1021 = n930 ^ n848 ;
  assign n928 = n844 & n877 ;
  assign n1022 = n1021 ^ n928 ;
  assign n1023 = n760 & ~n789 ;
  assign n1024 = n1023 ^ n846 ;
  assign n1029 = n1022 & n1024 ;
  assign n1030 = n1029 ^ n1024 ;
  assign n1031 = n1020 & n1030 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1034 = n1033 ^ n1032 ;
  assign n1035 = n1013 & n1034 ;
  assign n1040 = n1039 ^ n1035 ;
  assign n1041 = n998 & n1040 ;
  assign n1052 = n1051 ^ n1041 ;
  assign n1025 = n1024 ^ n1022 ;
  assign n1026 = ~n1020 & ~n1025 ;
  assign n1027 = n1013 & n1026 ;
  assign n1028 = n998 & n1027 ;
  assign n1053 = n1052 ^ n1028 ;
  assign n1145 = n970 & ~n1053 ;
  assign n1144 = n973 & n1053 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1055 = n973 & ~n1053 ;
  assign n1054 = n970 & n1053 ;
  assign n1056 = n1055 ^ n1054 ;
  assign n879 = n795 & ~n877 ;
  assign n878 = n792 & n877 ;
  assign n880 = n879 ^ n878 ;
  assign n615 = n531 & ~n613 ;
  assign n614 = n528 & n613 ;
  assign n616 = n615 ^ n614 ;
  assign n285 = x32 & ~n283 ;
  assign n284 = n221 & n283 ;
  assign n286 = n285 ^ n284 ;
  assign n344 = ~x40 & n286 ;
  assign n287 = n286 ^ x40 ;
  assign n289 = x33 & ~n283 ;
  assign n288 = n225 & n283 ;
  assign n290 = n289 ^ n288 ;
  assign n342 = ~x41 & n290 ;
  assign n343 = ~n287 & n342 ;
  assign n345 = n344 ^ n343 ;
  assign n291 = n290 ^ x41 ;
  assign n292 = ~n287 & ~n291 ;
  assign n294 = x34 & ~n283 ;
  assign n293 = n230 & n283 ;
  assign n295 = n294 ^ n293 ;
  assign n339 = ~x42 & n295 ;
  assign n296 = n295 ^ x42 ;
  assign n298 = x35 & ~n283 ;
  assign n297 = n234 & n283 ;
  assign n299 = n298 ^ n297 ;
  assign n337 = ~x43 & n299 ;
  assign n338 = ~n296 & n337 ;
  assign n340 = n339 ^ n338 ;
  assign n341 = n292 & n340 ;
  assign n346 = n345 ^ n341 ;
  assign n300 = n299 ^ x43 ;
  assign n301 = ~n296 & ~n300 ;
  assign n302 = n292 & n301 ;
  assign n304 = x36 & ~n283 ;
  assign n303 = n240 & n283 ;
  assign n305 = n304 ^ n303 ;
  assign n333 = ~x44 & n305 ;
  assign n306 = n305 ^ x44 ;
  assign n308 = x37 & ~n283 ;
  assign n307 = n244 & n283 ;
  assign n309 = n308 ^ n307 ;
  assign n331 = ~x45 & n309 ;
  assign n332 = ~n306 & n331 ;
  assign n334 = n333 ^ n332 ;
  assign n310 = n309 ^ x45 ;
  assign n311 = ~n306 & ~n310 ;
  assign n313 = x38 & ~n283 ;
  assign n312 = n249 & n283 ;
  assign n314 = n313 ^ n312 ;
  assign n328 = ~x46 & n314 ;
  assign n315 = n314 ^ x46 ;
  assign n317 = n316 ^ x39 ;
  assign n319 = n318 ^ n317 ;
  assign n324 = x47 & n319 ;
  assign n325 = n324 ^ n319 ;
  assign n326 = n315 & n325 ;
  assign n327 = n326 ^ n325 ;
  assign n329 = n328 ^ n327 ;
  assign n330 = n311 & n329 ;
  assign n335 = n334 ^ n330 ;
  assign n336 = n302 & n335 ;
  assign n347 = n346 ^ n336 ;
  assign n320 = n319 ^ x47 ;
  assign n321 = ~n315 & ~n320 ;
  assign n322 = n311 & n321 ;
  assign n323 = n302 & n322 ;
  assign n348 = n347 ^ n323 ;
  assign n350 = n286 & ~n348 ;
  assign n349 = x40 & n348 ;
  assign n351 = n350 ^ n349 ;
  assign n696 = ~n351 & n616 ;
  assign n617 = n616 ^ n351 ;
  assign n619 = n535 & ~n613 ;
  assign n618 = n538 & n613 ;
  assign n620 = n619 ^ n618 ;
  assign n622 = n290 & ~n348 ;
  assign n621 = x41 & n348 ;
  assign n623 = n622 ^ n621 ;
  assign n694 = n620 & ~n623 ;
  assign n695 = ~n617 & n694 ;
  assign n697 = n696 ^ n695 ;
  assign n624 = n623 ^ n620 ;
  assign n625 = ~n617 & ~n624 ;
  assign n627 = n546 & ~n613 ;
  assign n626 = n543 & n613 ;
  assign n628 = n627 ^ n626 ;
  assign n630 = n295 & ~n348 ;
  assign n629 = x42 & n348 ;
  assign n631 = n630 ^ n629 ;
  assign n691 = n628 & ~n631 ;
  assign n632 = n631 ^ n628 ;
  assign n634 = n553 & ~n613 ;
  assign n633 = n550 & n613 ;
  assign n635 = n634 ^ n633 ;
  assign n637 = n299 & ~n348 ;
  assign n636 = x43 & n348 ;
  assign n638 = n637 ^ n636 ;
  assign n689 = n635 & ~n638 ;
  assign n690 = ~n632 & n689 ;
  assign n692 = n691 ^ n690 ;
  assign n693 = n625 & n692 ;
  assign n698 = n697 ^ n693 ;
  assign n639 = n638 ^ n635 ;
  assign n640 = ~n632 & ~n639 ;
  assign n641 = n625 & n640 ;
  assign n643 = n562 & ~n613 ;
  assign n642 = n559 & n613 ;
  assign n644 = n643 ^ n642 ;
  assign n646 = n305 & ~n348 ;
  assign n645 = x44 & n348 ;
  assign n647 = n646 ^ n645 ;
  assign n685 = n644 & ~n647 ;
  assign n648 = n647 ^ n644 ;
  assign n650 = n569 & ~n613 ;
  assign n649 = n566 & n613 ;
  assign n651 = n650 ^ n649 ;
  assign n653 = n309 & ~n348 ;
  assign n652 = x45 & n348 ;
  assign n654 = n653 ^ n652 ;
  assign n683 = n651 & ~n654 ;
  assign n684 = ~n648 & n683 ;
  assign n686 = n685 ^ n684 ;
  assign n655 = n654 ^ n651 ;
  assign n656 = ~n648 & ~n655 ;
  assign n658 = n577 & ~n613 ;
  assign n657 = n574 & n613 ;
  assign n659 = n658 ^ n657 ;
  assign n661 = n314 & ~n348 ;
  assign n660 = x46 & n348 ;
  assign n662 = n661 ^ n660 ;
  assign n680 = n659 & ~n662 ;
  assign n663 = n662 ^ n659 ;
  assign n665 = n664 ^ n580 ;
  assign n667 = n666 ^ n665 ;
  assign n669 = n319 & n348 ;
  assign n670 = n669 ^ n319 ;
  assign n668 = x47 & n348 ;
  assign n671 = n670 ^ n668 ;
  assign n676 = n667 & n671 ;
  assign n677 = n676 ^ n667 ;
  assign n678 = n663 & n677 ;
  assign n679 = n678 ^ n677 ;
  assign n681 = n680 ^ n679 ;
  assign n682 = n656 & n681 ;
  assign n687 = n686 ^ n682 ;
  assign n688 = n641 & n687 ;
  assign n699 = n698 ^ n688 ;
  assign n672 = n671 ^ n667 ;
  assign n673 = ~n663 & ~n672 ;
  assign n674 = n656 & n673 ;
  assign n675 = n641 & n674 ;
  assign n700 = n699 ^ n675 ;
  assign n702 = n616 & ~n700 ;
  assign n701 = n351 & n700 ;
  assign n703 = n702 ^ n701 ;
  assign n960 = ~n703 & n880 ;
  assign n881 = n880 ^ n703 ;
  assign n883 = n799 & ~n877 ;
  assign n882 = n802 & n877 ;
  assign n884 = n883 ^ n882 ;
  assign n886 = n620 & ~n700 ;
  assign n885 = n623 & n700 ;
  assign n887 = n886 ^ n885 ;
  assign n958 = n884 & ~n887 ;
  assign n959 = ~n881 & n958 ;
  assign n961 = n960 ^ n959 ;
  assign n888 = n887 ^ n884 ;
  assign n889 = ~n881 & ~n888 ;
  assign n891 = n810 & ~n877 ;
  assign n890 = n807 & n877 ;
  assign n892 = n891 ^ n890 ;
  assign n894 = n628 & ~n700 ;
  assign n893 = n631 & n700 ;
  assign n895 = n894 ^ n893 ;
  assign n955 = n892 & ~n895 ;
  assign n896 = n895 ^ n892 ;
  assign n898 = n817 & ~n877 ;
  assign n897 = n814 & n877 ;
  assign n899 = n898 ^ n897 ;
  assign n901 = n635 & ~n700 ;
  assign n900 = n638 & n700 ;
  assign n902 = n901 ^ n900 ;
  assign n953 = n899 & ~n902 ;
  assign n954 = ~n896 & n953 ;
  assign n956 = n955 ^ n954 ;
  assign n957 = n889 & n956 ;
  assign n962 = n961 ^ n957 ;
  assign n903 = n902 ^ n899 ;
  assign n904 = ~n896 & ~n903 ;
  assign n905 = n889 & n904 ;
  assign n907 = n826 & ~n877 ;
  assign n906 = n823 & n877 ;
  assign n908 = n907 ^ n906 ;
  assign n910 = n644 & ~n700 ;
  assign n909 = n647 & n700 ;
  assign n911 = n910 ^ n909 ;
  assign n949 = n908 & ~n911 ;
  assign n912 = n911 ^ n908 ;
  assign n914 = n833 & ~n877 ;
  assign n913 = n830 & n877 ;
  assign n915 = n914 ^ n913 ;
  assign n917 = n651 & ~n700 ;
  assign n916 = n654 & n700 ;
  assign n918 = n917 ^ n916 ;
  assign n947 = n915 & ~n918 ;
  assign n948 = ~n912 & n947 ;
  assign n950 = n949 ^ n948 ;
  assign n919 = n918 ^ n915 ;
  assign n920 = ~n912 & ~n919 ;
  assign n922 = n841 & ~n877 ;
  assign n921 = n838 & n877 ;
  assign n923 = n922 ^ n921 ;
  assign n925 = n659 & ~n700 ;
  assign n924 = n662 & n700 ;
  assign n926 = n925 ^ n924 ;
  assign n944 = n923 & ~n926 ;
  assign n927 = n926 ^ n923 ;
  assign n929 = n928 ^ n844 ;
  assign n931 = n930 ^ n929 ;
  assign n933 = n667 & n700 ;
  assign n934 = n933 ^ n667 ;
  assign n932 = n671 & n700 ;
  assign n935 = n934 ^ n932 ;
  assign n940 = n931 & n935 ;
  assign n941 = n940 ^ n931 ;
  assign n942 = n927 & n941 ;
  assign n943 = n942 ^ n941 ;
  assign n945 = n944 ^ n943 ;
  assign n946 = n920 & n945 ;
  assign n951 = n950 ^ n946 ;
  assign n952 = n905 & n951 ;
  assign n963 = n962 ^ n952 ;
  assign n936 = n935 ^ n931 ;
  assign n937 = ~n927 & ~n936 ;
  assign n938 = n920 & n937 ;
  assign n939 = n905 & n938 ;
  assign n964 = n963 ^ n939 ;
  assign n966 = n880 & ~n964 ;
  assign n965 = n703 & n964 ;
  assign n967 = n966 ^ n965 ;
  assign n1136 = ~n967 & n1056 ;
  assign n1057 = n1056 ^ n967 ;
  assign n1059 = n977 & ~n1053 ;
  assign n1058 = n980 & n1053 ;
  assign n1060 = n1059 ^ n1058 ;
  assign n1062 = n884 & ~n964 ;
  assign n1061 = n887 & n964 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1134 = n1060 & ~n1063 ;
  assign n1135 = ~n1057 & n1134 ;
  assign n1137 = n1136 ^ n1135 ;
  assign n1064 = n1063 ^ n1060 ;
  assign n1065 = ~n1057 & ~n1064 ;
  assign n1067 = n988 & ~n1053 ;
  assign n1066 = n985 & n1053 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n1070 = n892 & ~n964 ;
  assign n1069 = n895 & n964 ;
  assign n1071 = n1070 ^ n1069 ;
  assign n1131 = n1068 & ~n1071 ;
  assign n1072 = n1071 ^ n1068 ;
  assign n1074 = n995 & ~n1053 ;
  assign n1073 = n992 & n1053 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1077 = n899 & ~n964 ;
  assign n1076 = n902 & n964 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1129 = n1075 & ~n1078 ;
  assign n1130 = ~n1072 & n1129 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1133 = n1065 & n1132 ;
  assign n1138 = n1137 ^ n1133 ;
  assign n1079 = n1078 ^ n1075 ;
  assign n1080 = ~n1072 & ~n1079 ;
  assign n1081 = n1065 & n1080 ;
  assign n1083 = n1004 & ~n1053 ;
  assign n1082 = n1001 & n1053 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1086 = n908 & ~n964 ;
  assign n1085 = n911 & n964 ;
  assign n1087 = n1086 ^ n1085 ;
  assign n1125 = n1084 & ~n1087 ;
  assign n1088 = n1087 ^ n1084 ;
  assign n1090 = n1011 & ~n1053 ;
  assign n1089 = n1008 & n1053 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1093 = n915 & ~n964 ;
  assign n1092 = n918 & n964 ;
  assign n1094 = n1093 ^ n1092 ;
  assign n1123 = n1091 & ~n1094 ;
  assign n1124 = ~n1088 & n1123 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1095 = n1094 ^ n1091 ;
  assign n1096 = ~n1088 & ~n1095 ;
  assign n1098 = n1019 & ~n1053 ;
  assign n1097 = n1016 & n1053 ;
  assign n1099 = n1098 ^ n1097 ;
  assign n1101 = n923 & ~n964 ;
  assign n1100 = n926 & n964 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1120 = n1099 & ~n1102 ;
  assign n1103 = n1102 ^ n1099 ;
  assign n1105 = n1022 & n1053 ;
  assign n1106 = n1105 ^ n1022 ;
  assign n1104 = n1024 & n1053 ;
  assign n1107 = n1106 ^ n1104 ;
  assign n1109 = n931 & n964 ;
  assign n1110 = n1109 ^ n931 ;
  assign n1108 = n935 & n964 ;
  assign n1111 = n1110 ^ n1108 ;
  assign n1116 = n1107 & n1111 ;
  assign n1117 = n1116 ^ n1107 ;
  assign n1118 = n1103 & n1117 ;
  assign n1119 = n1118 ^ n1117 ;
  assign n1121 = n1120 ^ n1119 ;
  assign n1122 = n1096 & n1121 ;
  assign n1127 = n1126 ^ n1122 ;
  assign n1128 = n1081 & n1127 ;
  assign n1139 = n1138 ^ n1128 ;
  assign n1112 = n1111 ^ n1107 ;
  assign n1113 = ~n1103 & ~n1112 ;
  assign n1114 = n1096 & n1113 ;
  assign n1115 = n1081 & n1114 ;
  assign n1140 = n1139 ^ n1115 ;
  assign n1142 = n1056 & ~n1140 ;
  assign n1141 = n967 & n1140 ;
  assign n1143 = n1142 ^ n1141 ;
  assign n1224 = ~n1143 & n1146 ;
  assign n1147 = n1146 ^ n1143 ;
  assign n1149 = n980 & ~n1053 ;
  assign n1148 = n977 & n1053 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1152 = n1060 & ~n1140 ;
  assign n1151 = n1063 & n1140 ;
  assign n1153 = n1152 ^ n1151 ;
  assign n1222 = n1150 & ~n1153 ;
  assign n1223 = ~n1147 & n1222 ;
  assign n1225 = n1224 ^ n1223 ;
  assign n1154 = n1153 ^ n1150 ;
  assign n1155 = ~n1147 & ~n1154 ;
  assign n1157 = n985 & ~n1053 ;
  assign n1156 = n988 & n1053 ;
  assign n1158 = n1157 ^ n1156 ;
  assign n1160 = n1068 & ~n1140 ;
  assign n1159 = n1071 & n1140 ;
  assign n1161 = n1160 ^ n1159 ;
  assign n1219 = n1158 & ~n1161 ;
  assign n1162 = n1161 ^ n1158 ;
  assign n1164 = n992 & ~n1053 ;
  assign n1163 = n995 & n1053 ;
  assign n1165 = n1164 ^ n1163 ;
  assign n1167 = n1075 & ~n1140 ;
  assign n1166 = n1078 & n1140 ;
  assign n1168 = n1167 ^ n1166 ;
  assign n1217 = n1165 & ~n1168 ;
  assign n1218 = ~n1162 & n1217 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1221 = n1155 & n1220 ;
  assign n1226 = n1225 ^ n1221 ;
  assign n1169 = n1168 ^ n1165 ;
  assign n1170 = ~n1162 & ~n1169 ;
  assign n1171 = n1155 & n1170 ;
  assign n1173 = n1001 & ~n1053 ;
  assign n1172 = n1004 & n1053 ;
  assign n1174 = n1173 ^ n1172 ;
  assign n1176 = n1084 & ~n1140 ;
  assign n1175 = n1087 & n1140 ;
  assign n1177 = n1176 ^ n1175 ;
  assign n1213 = n1174 & ~n1177 ;
  assign n1178 = n1177 ^ n1174 ;
  assign n1180 = n1008 & ~n1053 ;
  assign n1179 = n1011 & n1053 ;
  assign n1181 = n1180 ^ n1179 ;
  assign n1183 = n1091 & ~n1140 ;
  assign n1182 = n1094 & n1140 ;
  assign n1184 = n1183 ^ n1182 ;
  assign n1211 = n1181 & ~n1184 ;
  assign n1212 = ~n1178 & n1211 ;
  assign n1214 = n1213 ^ n1212 ;
  assign n1185 = n1184 ^ n1181 ;
  assign n1186 = ~n1178 & ~n1185 ;
  assign n1188 = n1016 & ~n1053 ;
  assign n1187 = n1019 & n1053 ;
  assign n1189 = n1188 ^ n1187 ;
  assign n1191 = n1099 & ~n1140 ;
  assign n1190 = n1102 & n1140 ;
  assign n1192 = n1191 ^ n1190 ;
  assign n1208 = n1189 & ~n1192 ;
  assign n1193 = n1192 ^ n1189 ;
  assign n1194 = n1024 & ~n1053 ;
  assign n1195 = n1194 ^ n1105 ;
  assign n1197 = n1107 & n1140 ;
  assign n1198 = n1197 ^ n1107 ;
  assign n1196 = n1111 & n1140 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1204 = n1195 & n1199 ;
  assign n1205 = n1204 ^ n1195 ;
  assign n1206 = n1193 & n1205 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1210 = n1186 & n1209 ;
  assign n1215 = n1214 ^ n1210 ;
  assign n1216 = n1171 & n1215 ;
  assign n1227 = n1226 ^ n1216 ;
  assign n1200 = n1199 ^ n1195 ;
  assign n1201 = ~n1193 & ~n1200 ;
  assign n1202 = n1186 & n1201 ;
  assign n1203 = n1171 & n1202 ;
  assign n1228 = n1227 ^ n1203 ;
  assign n1230 = n1146 & n1228 ;
  assign n1231 = n1230 ^ n1146 ;
  assign n1229 = n1143 & n1228 ;
  assign n1232 = n1231 ^ n1229 ;
  assign n1234 = n1150 & n1228 ;
  assign n1235 = n1234 ^ n1150 ;
  assign n1233 = n1153 & n1228 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1238 = n1158 & n1228 ;
  assign n1239 = n1238 ^ n1158 ;
  assign n1237 = n1161 & n1228 ;
  assign n1240 = n1239 ^ n1237 ;
  assign n1242 = n1165 & n1228 ;
  assign n1243 = n1242 ^ n1165 ;
  assign n1241 = n1168 & n1228 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1246 = n1174 & n1228 ;
  assign n1247 = n1246 ^ n1174 ;
  assign n1245 = n1177 & n1228 ;
  assign n1248 = n1247 ^ n1245 ;
  assign n1250 = n1181 & n1228 ;
  assign n1251 = n1250 ^ n1181 ;
  assign n1249 = n1184 & n1228 ;
  assign n1252 = n1251 ^ n1249 ;
  assign n1254 = n1189 & n1228 ;
  assign n1255 = n1254 ^ n1189 ;
  assign n1253 = n1192 & n1228 ;
  assign n1256 = n1255 ^ n1253 ;
  assign n1258 = n1195 & n1228 ;
  assign n1259 = n1258 ^ n1195 ;
  assign n1257 = n1199 & n1228 ;
  assign n1260 = n1259 ^ n1257 ;
  assign n1261 = n1229 ^ n1143 ;
  assign n1262 = n1261 ^ n1230 ;
  assign n1263 = n1233 ^ n1153 ;
  assign n1264 = n1263 ^ n1234 ;
  assign n1265 = n1237 ^ n1161 ;
  assign n1266 = n1265 ^ n1238 ;
  assign n1267 = n1241 ^ n1168 ;
  assign n1268 = n1267 ^ n1242 ;
  assign n1269 = n1245 ^ n1177 ;
  assign n1270 = n1269 ^ n1246 ;
  assign n1271 = n1249 ^ n1184 ;
  assign n1272 = n1271 ^ n1250 ;
  assign n1273 = n1253 ^ n1192 ;
  assign n1274 = n1273 ^ n1254 ;
  assign n1275 = n1257 ^ n1199 ;
  assign n1276 = n1275 ^ n1258 ;
  assign n1278 = n967 & ~n1140 ;
  assign n1277 = n1056 & n1140 ;
  assign n1279 = n1278 ^ n1277 ;
  assign n1281 = n1063 & ~n1140 ;
  assign n1280 = n1060 & n1140 ;
  assign n1282 = n1281 ^ n1280 ;
  assign n1284 = n1071 & ~n1140 ;
  assign n1283 = n1068 & n1140 ;
  assign n1285 = n1284 ^ n1283 ;
  assign n1287 = n1078 & ~n1140 ;
  assign n1286 = n1075 & n1140 ;
  assign n1288 = n1287 ^ n1286 ;
  assign n1290 = n1087 & ~n1140 ;
  assign n1289 = n1084 & n1140 ;
  assign n1291 = n1290 ^ n1289 ;
  assign n1293 = n1094 & ~n1140 ;
  assign n1292 = n1091 & n1140 ;
  assign n1294 = n1293 ^ n1292 ;
  assign n1296 = n1102 & ~n1140 ;
  assign n1295 = n1099 & n1140 ;
  assign n1297 = n1296 ^ n1295 ;
  assign n1298 = n1111 & ~n1140 ;
  assign n1299 = n1298 ^ n1197 ;
  assign n1301 = n703 & ~n964 ;
  assign n1300 = n880 & n964 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1304 = n887 & ~n964 ;
  assign n1303 = n884 & n964 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1307 = n895 & ~n964 ;
  assign n1306 = n892 & n964 ;
  assign n1308 = n1307 ^ n1306 ;
  assign n1310 = n902 & ~n964 ;
  assign n1309 = n899 & n964 ;
  assign n1311 = n1310 ^ n1309 ;
  assign n1313 = n911 & ~n964 ;
  assign n1312 = n908 & n964 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1316 = n918 & ~n964 ;
  assign n1315 = n915 & n964 ;
  assign n1317 = n1316 ^ n1315 ;
  assign n1319 = n926 & ~n964 ;
  assign n1318 = n923 & n964 ;
  assign n1320 = n1319 ^ n1318 ;
  assign n1321 = n935 & ~n964 ;
  assign n1322 = n1321 ^ n1109 ;
  assign n1324 = n351 & ~n700 ;
  assign n1323 = n616 & n700 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1327 = n623 & ~n700 ;
  assign n1326 = n620 & n700 ;
  assign n1328 = n1327 ^ n1326 ;
  assign n1330 = n631 & ~n700 ;
  assign n1329 = n628 & n700 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1333 = n638 & ~n700 ;
  assign n1332 = n635 & n700 ;
  assign n1334 = n1333 ^ n1332 ;
  assign n1336 = n647 & ~n700 ;
  assign n1335 = n644 & n700 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1339 = n654 & ~n700 ;
  assign n1338 = n651 & n700 ;
  assign n1340 = n1339 ^ n1338 ;
  assign n1342 = n662 & ~n700 ;
  assign n1341 = n659 & n700 ;
  assign n1343 = n1342 ^ n1341 ;
  assign n1344 = n671 & ~n700 ;
  assign n1345 = n1344 ^ n933 ;
  assign n1347 = x40 & ~n348 ;
  assign n1346 = n286 & n348 ;
  assign n1348 = n1347 ^ n1346 ;
  assign n1350 = x41 & ~n348 ;
  assign n1349 = n290 & n348 ;
  assign n1351 = n1350 ^ n1349 ;
  assign n1353 = x42 & ~n348 ;
  assign n1352 = n295 & n348 ;
  assign n1354 = n1353 ^ n1352 ;
  assign n1356 = x43 & ~n348 ;
  assign n1355 = n299 & n348 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1359 = x44 & ~n348 ;
  assign n1358 = n305 & n348 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1362 = x45 & ~n348 ;
  assign n1361 = n309 & n348 ;
  assign n1363 = n1362 ^ n1361 ;
  assign n1365 = x46 & ~n348 ;
  assign n1364 = n314 & n348 ;
  assign n1366 = n1365 ^ n1364 ;
  assign n1367 = x47 & ~n348 ;
  assign n1368 = n1367 ^ n669 ;
  assign y0 = n1232 ;
  assign y1 = n1236 ;
  assign y2 = n1240 ;
  assign y3 = n1244 ;
  assign y4 = n1248 ;
  assign y5 = n1252 ;
  assign y6 = n1256 ;
  assign y7 = n1260 ;
  assign y8 = n1262 ;
  assign y9 = n1264 ;
  assign y10 = n1266 ;
  assign y11 = n1268 ;
  assign y12 = n1270 ;
  assign y13 = n1272 ;
  assign y14 = n1274 ;
  assign y15 = n1276 ;
  assign y16 = n1279 ;
  assign y17 = n1282 ;
  assign y18 = n1285 ;
  assign y19 = n1288 ;
  assign y20 = n1291 ;
  assign y21 = n1294 ;
  assign y22 = n1297 ;
  assign y23 = n1299 ;
  assign y24 = n1302 ;
  assign y25 = n1305 ;
  assign y26 = n1308 ;
  assign y27 = n1311 ;
  assign y28 = n1314 ;
  assign y29 = n1317 ;
  assign y30 = n1320 ;
  assign y31 = n1322 ;
  assign y32 = n1325 ;
  assign y33 = n1328 ;
  assign y34 = n1331 ;
  assign y35 = n1334 ;
  assign y36 = n1337 ;
  assign y37 = n1340 ;
  assign y38 = n1343 ;
  assign y39 = n1345 ;
  assign y40 = n1348 ;
  assign y41 = n1351 ;
  assign y42 = n1354 ;
  assign y43 = n1357 ;
  assign y44 = n1360 ;
  assign y45 = n1363 ;
  assign y46 = n1366 ;
  assign y47 = n1368 ;
endmodule
