module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 ;
  assign n54 = x8 ^ x0 ;
  assign n55 = x9 ^ x1 ;
  assign n56 = ~n54 & ~n55 ;
  assign n49 = x10 ^ x2 ;
  assign n65 = x11 ^ x3 ;
  assign n66 = ~n49 & ~n65 ;
  assign n67 = n56 & n66 ;
  assign n85 = x4 & ~x12 ;
  assign n68 = x12 ^ x4 ;
  assign n83 = x5 & ~x13 ;
  assign n84 = ~n68 & n83 ;
  assign n86 = n85 ^ n84 ;
  assign n69 = x13 ^ x5 ;
  assign n70 = ~n68 & ~n69 ;
  assign n80 = x6 & ~x14 ;
  assign n71 = x14 ^ x6 ;
  assign n78 = x7 & ~x15 ;
  assign n79 = ~n71 & n78 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n70 & n81 ;
  assign n87 = n86 ^ n82 ;
  assign n675 = n67 & n87 ;
  assign n52 = x2 & ~x10 ;
  assign n50 = x3 & ~x11 ;
  assign n51 = ~n49 & n50 ;
  assign n53 = n52 ^ n51 ;
  assign n673 = n53 & n56 ;
  assign n61 = x0 & ~x8 ;
  assign n59 = x1 & ~x9 ;
  assign n60 = ~n54 & n59 ;
  assign n62 = n61 ^ n60 ;
  assign n674 = n673 ^ n62 ;
  assign n676 = n675 ^ n674 ;
  assign n72 = x15 ^ x7 ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = n70 & n73 ;
  assign n75 = n67 & n74 ;
  assign n677 = n676 ^ n75 ;
  assign n679 = x0 & ~n677 ;
  assign n678 = x8 & n677 ;
  assign n680 = n679 ^ n678 ;
  assign n97 = x8 & n67 ;
  assign n98 = n87 & n97 ;
  assign n95 = x8 & ~n75 ;
  assign n93 = x8 & n62 ;
  assign n91 = x8 & n56 ;
  assign n92 = n53 & n91 ;
  assign n94 = n93 ^ n92 ;
  assign n96 = n95 ^ n94 ;
  assign n99 = n98 ^ n96 ;
  assign n88 = x0 & n67 ;
  assign n89 = n87 & n88 ;
  assign n76 = x0 & ~n75 ;
  assign n63 = x0 & ~n62 ;
  assign n57 = x0 & n56 ;
  assign n58 = n53 & n57 ;
  assign n64 = n63 ^ n58 ;
  assign n77 = n76 ^ n64 ;
  assign n90 = n89 ^ n77 ;
  assign n100 = n99 ^ n90 ;
  assign n123 = ~x16 & n100 ;
  assign n101 = n100 ^ x16 ;
  assign n117 = x9 & n67 ;
  assign n118 = n87 & n117 ;
  assign n115 = x9 & ~n75 ;
  assign n113 = x9 & n62 ;
  assign n111 = x9 & n56 ;
  assign n112 = n53 & n111 ;
  assign n114 = n113 ^ n112 ;
  assign n116 = n115 ^ n114 ;
  assign n119 = n118 ^ n116 ;
  assign n108 = x1 & n67 ;
  assign n109 = n87 & n108 ;
  assign n106 = x1 & ~n75 ;
  assign n104 = x1 & ~n62 ;
  assign n102 = x1 & n56 ;
  assign n103 = n53 & n102 ;
  assign n105 = n104 ^ n103 ;
  assign n107 = n106 ^ n105 ;
  assign n110 = n109 ^ n107 ;
  assign n120 = n119 ^ n110 ;
  assign n121 = ~x17 & n120 ;
  assign n122 = ~n101 & n121 ;
  assign n124 = n123 ^ n122 ;
  assign n685 = n100 & n124 ;
  assign n141 = x10 & n67 ;
  assign n142 = n87 & n141 ;
  assign n139 = x10 & ~n75 ;
  assign n137 = x10 & n62 ;
  assign n135 = x10 & n56 ;
  assign n136 = n53 & n135 ;
  assign n138 = n137 ^ n136 ;
  assign n140 = n139 ^ n138 ;
  assign n143 = n142 ^ n140 ;
  assign n132 = x2 & n67 ;
  assign n133 = n87 & n132 ;
  assign n130 = x2 & ~n75 ;
  assign n128 = x2 & ~n62 ;
  assign n126 = x2 & n56 ;
  assign n127 = n53 & n126 ;
  assign n129 = n128 ^ n127 ;
  assign n131 = n130 ^ n129 ;
  assign n134 = n133 ^ n131 ;
  assign n144 = n143 ^ n134 ;
  assign n167 = ~x18 & n144 ;
  assign n145 = n144 ^ x18 ;
  assign n161 = x11 & n67 ;
  assign n162 = n87 & n161 ;
  assign n159 = x11 & ~n75 ;
  assign n157 = x11 & n62 ;
  assign n155 = x11 & n56 ;
  assign n156 = n53 & n155 ;
  assign n158 = n157 ^ n156 ;
  assign n160 = n159 ^ n158 ;
  assign n163 = n162 ^ n160 ;
  assign n152 = x3 & n67 ;
  assign n153 = n87 & n152 ;
  assign n150 = x3 & ~n75 ;
  assign n148 = x3 & ~n62 ;
  assign n146 = x3 & n56 ;
  assign n147 = n53 & n146 ;
  assign n149 = n148 ^ n147 ;
  assign n151 = n150 ^ n149 ;
  assign n154 = n153 ^ n151 ;
  assign n164 = n163 ^ n154 ;
  assign n165 = ~x19 & n164 ;
  assign n166 = ~n145 & n165 ;
  assign n168 = n167 ^ n166 ;
  assign n169 = n120 ^ x17 ;
  assign n170 = ~n101 & ~n169 ;
  assign n171 = n100 & n170 ;
  assign n172 = n168 & n171 ;
  assign n686 = n685 ^ n172 ;
  assign n174 = n164 ^ x19 ;
  assign n175 = ~n145 & ~n174 ;
  assign n176 = n170 & n175 ;
  assign n192 = x12 & n67 ;
  assign n193 = n87 & n192 ;
  assign n190 = x12 & ~n75 ;
  assign n188 = x12 & n62 ;
  assign n186 = x12 & n56 ;
  assign n187 = n53 & n186 ;
  assign n189 = n188 ^ n187 ;
  assign n191 = n190 ^ n189 ;
  assign n194 = n193 ^ n191 ;
  assign n183 = x4 & n67 ;
  assign n184 = n87 & n183 ;
  assign n181 = x4 & ~n75 ;
  assign n179 = x4 & ~n62 ;
  assign n177 = x4 & n56 ;
  assign n178 = n53 & n177 ;
  assign n180 = n179 ^ n178 ;
  assign n182 = n181 ^ n180 ;
  assign n185 = n184 ^ n182 ;
  assign n195 = n194 ^ n185 ;
  assign n196 = n195 ^ x20 ;
  assign n212 = x13 & n67 ;
  assign n213 = n87 & n212 ;
  assign n210 = x13 & ~n75 ;
  assign n208 = x13 & n62 ;
  assign n206 = x13 & n56 ;
  assign n207 = n53 & n206 ;
  assign n209 = n208 ^ n207 ;
  assign n211 = n210 ^ n209 ;
  assign n214 = n213 ^ n211 ;
  assign n203 = x5 & n67 ;
  assign n204 = n87 & n203 ;
  assign n201 = x5 & ~n75 ;
  assign n199 = x5 & ~n62 ;
  assign n197 = x5 & n56 ;
  assign n198 = n53 & n197 ;
  assign n200 = n199 ^ n198 ;
  assign n202 = n201 ^ n200 ;
  assign n205 = n204 ^ n202 ;
  assign n215 = n214 ^ n205 ;
  assign n216 = n215 ^ x21 ;
  assign n217 = ~n196 & ~n216 ;
  assign n233 = x14 & n67 ;
  assign n234 = n87 & n233 ;
  assign n231 = x14 & ~n75 ;
  assign n229 = x14 & n62 ;
  assign n227 = x14 & n56 ;
  assign n228 = n53 & n227 ;
  assign n230 = n229 ^ n228 ;
  assign n232 = n231 ^ n230 ;
  assign n235 = n234 ^ n232 ;
  assign n224 = x6 & n67 ;
  assign n225 = n87 & n224 ;
  assign n222 = x6 & ~n75 ;
  assign n220 = x6 & ~n62 ;
  assign n218 = x6 & n56 ;
  assign n219 = n53 & n218 ;
  assign n221 = n220 ^ n219 ;
  assign n223 = n222 ^ n221 ;
  assign n226 = n225 ^ n223 ;
  assign n236 = n235 ^ n226 ;
  assign n237 = n236 ^ x22 ;
  assign n253 = x15 & n67 ;
  assign n254 = n87 & n253 ;
  assign n251 = x15 & ~n75 ;
  assign n249 = x15 & n62 ;
  assign n247 = x15 & n56 ;
  assign n248 = n53 & n247 ;
  assign n250 = n249 ^ n248 ;
  assign n252 = n251 ^ n250 ;
  assign n255 = n254 ^ n252 ;
  assign n244 = x7 & n67 ;
  assign n245 = n87 & n244 ;
  assign n242 = x7 & ~n75 ;
  assign n240 = x7 & ~n62 ;
  assign n238 = x7 & n56 ;
  assign n239 = n53 & n238 ;
  assign n241 = n240 ^ n239 ;
  assign n243 = n242 ^ n241 ;
  assign n246 = n245 ^ n243 ;
  assign n256 = n255 ^ n246 ;
  assign n257 = n256 ^ x23 ;
  assign n258 = ~n237 & ~n257 ;
  assign n259 = n217 & n258 ;
  assign n260 = n176 & n259 ;
  assign n261 = n100 & ~n260 ;
  assign n687 = n686 ^ n261 ;
  assign n263 = n100 & n176 ;
  assign n271 = ~x20 & n195 ;
  assign n269 = ~x21 & n215 ;
  assign n270 = ~n196 & n269 ;
  assign n272 = n271 ^ n270 ;
  assign n266 = ~x22 & n236 ;
  assign n264 = ~x23 & n256 ;
  assign n265 = ~n237 & n264 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = n217 & n267 ;
  assign n273 = n272 ^ n268 ;
  assign n274 = n263 & n273 ;
  assign n688 = n687 ^ n274 ;
  assign n681 = x16 & ~n124 ;
  assign n277 = x16 & n170 ;
  assign n278 = n168 & n277 ;
  assign n682 = n681 ^ n278 ;
  assign n280 = x16 & ~n260 ;
  assign n683 = n682 ^ n280 ;
  assign n282 = x16 & n176 ;
  assign n283 = n273 & n282 ;
  assign n684 = n683 ^ n283 ;
  assign n689 = n688 ^ n684 ;
  assign n868 = n680 & ~n689 ;
  assign n690 = n689 ^ n680 ;
  assign n695 = n120 & n124 ;
  assign n288 = n120 & n170 ;
  assign n289 = n168 & n288 ;
  assign n696 = n695 ^ n289 ;
  assign n291 = n120 & ~n260 ;
  assign n697 = n696 ^ n291 ;
  assign n293 = n120 & n176 ;
  assign n294 = n273 & n293 ;
  assign n698 = n697 ^ n294 ;
  assign n691 = x17 & ~n124 ;
  assign n297 = x17 & n170 ;
  assign n298 = n168 & n297 ;
  assign n692 = n691 ^ n298 ;
  assign n300 = x17 & ~n260 ;
  assign n693 = n692 ^ n300 ;
  assign n302 = x17 & n176 ;
  assign n303 = n273 & n302 ;
  assign n694 = n693 ^ n303 ;
  assign n699 = n698 ^ n694 ;
  assign n701 = x1 & ~n677 ;
  assign n700 = x9 & n677 ;
  assign n702 = n701 ^ n700 ;
  assign n866 = ~n699 & n702 ;
  assign n867 = ~n690 & n866 ;
  assign n869 = n868 ^ n867 ;
  assign n703 = n702 ^ n699 ;
  assign n704 = ~n690 & ~n703 ;
  assign n706 = x2 & ~n677 ;
  assign n705 = x10 & n677 ;
  assign n707 = n706 ^ n705 ;
  assign n712 = n124 & n144 ;
  assign n309 = n144 & n170 ;
  assign n310 = n168 & n309 ;
  assign n713 = n712 ^ n310 ;
  assign n312 = n144 & ~n260 ;
  assign n714 = n713 ^ n312 ;
  assign n314 = n144 & n176 ;
  assign n315 = n273 & n314 ;
  assign n715 = n714 ^ n315 ;
  assign n708 = x18 & ~n124 ;
  assign n318 = x18 & n170 ;
  assign n319 = n168 & n318 ;
  assign n709 = n708 ^ n319 ;
  assign n321 = x18 & ~n260 ;
  assign n710 = n709 ^ n321 ;
  assign n323 = x18 & n176 ;
  assign n324 = n273 & n323 ;
  assign n711 = n710 ^ n324 ;
  assign n716 = n715 ^ n711 ;
  assign n863 = n707 & ~n716 ;
  assign n717 = n716 ^ n707 ;
  assign n719 = x3 & ~n677 ;
  assign n718 = x11 & n677 ;
  assign n720 = n719 ^ n718 ;
  assign n725 = n124 & n164 ;
  assign n329 = n164 & n170 ;
  assign n330 = n168 & n329 ;
  assign n726 = n725 ^ n330 ;
  assign n332 = n164 & ~n260 ;
  assign n727 = n726 ^ n332 ;
  assign n334 = n164 & n176 ;
  assign n335 = n273 & n334 ;
  assign n728 = n727 ^ n335 ;
  assign n721 = x19 & ~n124 ;
  assign n338 = x19 & n170 ;
  assign n339 = n168 & n338 ;
  assign n722 = n721 ^ n339 ;
  assign n341 = x19 & ~n260 ;
  assign n723 = n722 ^ n341 ;
  assign n343 = x19 & n176 ;
  assign n344 = n273 & n343 ;
  assign n724 = n723 ^ n344 ;
  assign n729 = n728 ^ n724 ;
  assign n861 = n720 & ~n729 ;
  assign n862 = ~n717 & n861 ;
  assign n864 = n863 ^ n862 ;
  assign n865 = n704 & n864 ;
  assign n870 = n869 ^ n865 ;
  assign n730 = n729 ^ n720 ;
  assign n731 = ~n717 & ~n730 ;
  assign n732 = n704 & n731 ;
  assign n734 = x4 & ~n677 ;
  assign n733 = x12 & n677 ;
  assign n735 = n734 ^ n733 ;
  assign n740 = n124 & n195 ;
  assign n351 = n170 & n195 ;
  assign n352 = n168 & n351 ;
  assign n741 = n740 ^ n352 ;
  assign n354 = n195 & ~n260 ;
  assign n742 = n741 ^ n354 ;
  assign n356 = n176 & n195 ;
  assign n357 = n273 & n356 ;
  assign n743 = n742 ^ n357 ;
  assign n736 = x20 & ~n124 ;
  assign n360 = x20 & n170 ;
  assign n361 = n168 & n360 ;
  assign n737 = n736 ^ n361 ;
  assign n363 = x20 & ~n260 ;
  assign n738 = n737 ^ n363 ;
  assign n365 = x20 & n176 ;
  assign n366 = n273 & n365 ;
  assign n739 = n738 ^ n366 ;
  assign n744 = n743 ^ n739 ;
  assign n857 = n735 & ~n744 ;
  assign n745 = n744 ^ n735 ;
  assign n747 = x5 & ~n677 ;
  assign n746 = x13 & n677 ;
  assign n748 = n747 ^ n746 ;
  assign n753 = n124 & n215 ;
  assign n371 = n170 & n215 ;
  assign n372 = n168 & n371 ;
  assign n754 = n753 ^ n372 ;
  assign n374 = n215 & ~n260 ;
  assign n755 = n754 ^ n374 ;
  assign n376 = n176 & n215 ;
  assign n377 = n273 & n376 ;
  assign n756 = n755 ^ n377 ;
  assign n749 = x21 & ~n124 ;
  assign n380 = x21 & n170 ;
  assign n381 = n168 & n380 ;
  assign n750 = n749 ^ n381 ;
  assign n383 = x21 & ~n260 ;
  assign n751 = n750 ^ n383 ;
  assign n385 = x21 & n176 ;
  assign n386 = n273 & n385 ;
  assign n752 = n751 ^ n386 ;
  assign n757 = n756 ^ n752 ;
  assign n855 = n748 & ~n757 ;
  assign n856 = ~n745 & n855 ;
  assign n858 = n857 ^ n856 ;
  assign n758 = n757 ^ n748 ;
  assign n759 = ~n745 & ~n758 ;
  assign n770 = x6 & ~n677 ;
  assign n769 = x14 & n677 ;
  assign n771 = n770 ^ n769 ;
  assign n846 = ~n236 & n771 ;
  assign n850 = n176 & n846 ;
  assign n851 = n273 & n850 ;
  assign n436 = n168 & n170 ;
  assign n437 = n436 ^ n124 ;
  assign n848 = ~n437 & n846 ;
  assign n847 = n260 & n846 ;
  assign n849 = n848 ^ n847 ;
  assign n852 = n851 ^ n849 ;
  assign n786 = x7 & ~n674 ;
  assign n785 = x7 & n75 ;
  assign n787 = n786 ^ n785 ;
  assign n788 = n787 ^ n245 ;
  assign n782 = x15 & ~n674 ;
  assign n783 = n782 ^ n251 ;
  assign n784 = n783 ^ n254 ;
  assign n789 = n788 ^ n784 ;
  assign n811 = ~n256 & n789 ;
  assign n818 = n176 & n811 ;
  assign n819 = n273 & n818 ;
  assign n816 = ~n260 & n811 ;
  assign n814 = n124 & n811 ;
  assign n812 = n170 & n811 ;
  assign n813 = n168 & n812 ;
  assign n815 = n814 ^ n813 ;
  assign n817 = n816 ^ n815 ;
  assign n820 = n819 ^ n817 ;
  assign n801 = ~x23 & n789 ;
  assign n808 = n176 & n801 ;
  assign n809 = n273 & n808 ;
  assign n806 = ~n260 & n801 ;
  assign n804 = ~n124 & n801 ;
  assign n802 = n170 & n801 ;
  assign n803 = n168 & n802 ;
  assign n805 = n804 ^ n803 ;
  assign n807 = n806 ^ n805 ;
  assign n810 = n809 ^ n807 ;
  assign n821 = n820 ^ n810 ;
  assign n843 = n771 & n821 ;
  assign n838 = n176 & ~n236 ;
  assign n839 = n273 & n838 ;
  assign n836 = ~n236 & ~n260 ;
  assign n834 = n124 & ~n236 ;
  assign n832 = n170 & ~n236 ;
  assign n833 = n168 & n832 ;
  assign n835 = n834 ^ n833 ;
  assign n837 = n836 ^ n835 ;
  assign n840 = n839 ^ n837 ;
  assign n841 = n821 & n840 ;
  assign n828 = ~x22 & n176 ;
  assign n829 = n273 & n828 ;
  assign n826 = ~x22 & ~n260 ;
  assign n824 = ~x22 & ~n124 ;
  assign n822 = ~x22 & n170 ;
  assign n823 = n168 & n822 ;
  assign n825 = n824 ^ n823 ;
  assign n827 = n826 ^ n825 ;
  assign n830 = n829 ^ n827 ;
  assign n831 = n821 & n830 ;
  assign n842 = n841 ^ n831 ;
  assign n844 = n843 ^ n842 ;
  assign n794 = ~x22 & n771 ;
  assign n798 = n176 & n794 ;
  assign n799 = n273 & n798 ;
  assign n796 = ~n260 & n794 ;
  assign n795 = ~n437 & n794 ;
  assign n797 = n796 ^ n795 ;
  assign n800 = n799 ^ n797 ;
  assign n845 = n844 ^ n800 ;
  assign n853 = n852 ^ n845 ;
  assign n854 = n759 & n853 ;
  assign n859 = n858 ^ n854 ;
  assign n860 = n732 & n859 ;
  assign n871 = n870 ^ n860 ;
  assign n764 = n124 & n236 ;
  assign n392 = n170 & n236 ;
  assign n393 = n168 & n392 ;
  assign n765 = n764 ^ n393 ;
  assign n395 = n236 & ~n260 ;
  assign n766 = n765 ^ n395 ;
  assign n397 = n176 & n236 ;
  assign n398 = n273 & n397 ;
  assign n767 = n766 ^ n398 ;
  assign n760 = x22 & ~n124 ;
  assign n401 = x22 & n170 ;
  assign n402 = n168 & n401 ;
  assign n761 = n760 ^ n402 ;
  assign n404 = x22 & ~n260 ;
  assign n762 = n761 ^ n404 ;
  assign n406 = x22 & n176 ;
  assign n407 = n273 & n406 ;
  assign n763 = n762 ^ n407 ;
  assign n768 = n767 ^ n763 ;
  assign n772 = n771 ^ n768 ;
  assign n777 = n124 & n256 ;
  assign n412 = n170 & n256 ;
  assign n413 = n168 & n412 ;
  assign n778 = n777 ^ n413 ;
  assign n415 = n256 & ~n260 ;
  assign n779 = n778 ^ n415 ;
  assign n417 = n176 & n256 ;
  assign n418 = n273 & n417 ;
  assign n780 = n779 ^ n418 ;
  assign n773 = x23 & ~n124 ;
  assign n421 = x23 & n170 ;
  assign n422 = n168 & n421 ;
  assign n774 = n773 ^ n422 ;
  assign n424 = x23 & ~n260 ;
  assign n775 = n774 ^ n424 ;
  assign n426 = x23 & n176 ;
  assign n427 = n273 & n426 ;
  assign n776 = n775 ^ n427 ;
  assign n781 = n780 ^ n776 ;
  assign n790 = n789 ^ n781 ;
  assign n791 = ~n772 & ~n790 ;
  assign n792 = n759 & n791 ;
  assign n793 = n732 & n792 ;
  assign n872 = n871 ^ n793 ;
  assign n1398 = n680 & ~n872 ;
  assign n1397 = n689 & n872 ;
  assign n1399 = n1398 ^ n1397 ;
  assign n874 = n689 & ~n872 ;
  assign n873 = n680 & n872 ;
  assign n875 = n874 ^ n873 ;
  assign n276 = x16 & n124 ;
  assign n279 = n278 ^ n276 ;
  assign n281 = n280 ^ n279 ;
  assign n284 = n283 ^ n281 ;
  assign n125 = n100 & ~n124 ;
  assign n173 = n172 ^ n125 ;
  assign n262 = n261 ^ n173 ;
  assign n275 = n274 ^ n262 ;
  assign n285 = n284 ^ n275 ;
  assign n492 = ~x24 & n285 ;
  assign n286 = n285 ^ x24 ;
  assign n296 = x17 & n124 ;
  assign n299 = n298 ^ n296 ;
  assign n301 = n300 ^ n299 ;
  assign n304 = n303 ^ n301 ;
  assign n287 = n120 & ~n124 ;
  assign n290 = n289 ^ n287 ;
  assign n292 = n291 ^ n290 ;
  assign n295 = n294 ^ n292 ;
  assign n305 = n304 ^ n295 ;
  assign n490 = ~x25 & n305 ;
  assign n491 = ~n286 & n490 ;
  assign n493 = n492 ^ n491 ;
  assign n306 = n305 ^ x25 ;
  assign n307 = ~n286 & ~n306 ;
  assign n317 = x18 & n124 ;
  assign n320 = n319 ^ n317 ;
  assign n322 = n321 ^ n320 ;
  assign n325 = n324 ^ n322 ;
  assign n308 = ~n124 & n144 ;
  assign n311 = n310 ^ n308 ;
  assign n313 = n312 ^ n311 ;
  assign n316 = n315 ^ n313 ;
  assign n326 = n325 ^ n316 ;
  assign n487 = ~x26 & n326 ;
  assign n327 = n326 ^ x26 ;
  assign n337 = x19 & n124 ;
  assign n340 = n339 ^ n337 ;
  assign n342 = n341 ^ n340 ;
  assign n345 = n344 ^ n342 ;
  assign n328 = ~n124 & n164 ;
  assign n331 = n330 ^ n328 ;
  assign n333 = n332 ^ n331 ;
  assign n336 = n335 ^ n333 ;
  assign n346 = n345 ^ n336 ;
  assign n485 = ~x27 & n346 ;
  assign n486 = ~n327 & n485 ;
  assign n488 = n487 ^ n486 ;
  assign n489 = n307 & n488 ;
  assign n494 = n493 ^ n489 ;
  assign n347 = n346 ^ x27 ;
  assign n348 = ~n327 & ~n347 ;
  assign n349 = n307 & n348 ;
  assign n359 = x20 & n124 ;
  assign n362 = n361 ^ n359 ;
  assign n364 = n363 ^ n362 ;
  assign n367 = n366 ^ n364 ;
  assign n350 = ~n124 & n195 ;
  assign n353 = n352 ^ n350 ;
  assign n355 = n354 ^ n353 ;
  assign n358 = n357 ^ n355 ;
  assign n368 = n367 ^ n358 ;
  assign n481 = ~x28 & n368 ;
  assign n369 = n368 ^ x28 ;
  assign n379 = x21 & n124 ;
  assign n382 = n381 ^ n379 ;
  assign n384 = n383 ^ n382 ;
  assign n387 = n386 ^ n384 ;
  assign n370 = ~n124 & n215 ;
  assign n373 = n372 ^ n370 ;
  assign n375 = n374 ^ n373 ;
  assign n378 = n377 ^ n375 ;
  assign n388 = n387 ^ n378 ;
  assign n479 = ~x29 & n388 ;
  assign n480 = ~n369 & n479 ;
  assign n482 = n481 ^ n480 ;
  assign n389 = n388 ^ x29 ;
  assign n390 = ~n369 & ~n389 ;
  assign n470 = ~x30 & n236 ;
  assign n474 = n176 & n470 ;
  assign n475 = n273 & n474 ;
  assign n472 = ~n260 & n470 ;
  assign n471 = ~n437 & n470 ;
  assign n473 = n472 ^ n471 ;
  assign n476 = n475 ^ n473 ;
  assign n453 = ~x31 & n256 ;
  assign n460 = n176 & n453 ;
  assign n461 = n273 & n460 ;
  assign n458 = ~n260 & n453 ;
  assign n456 = ~n124 & n453 ;
  assign n454 = n170 & n453 ;
  assign n455 = n168 & n454 ;
  assign n457 = n456 ^ n455 ;
  assign n459 = n458 ^ n457 ;
  assign n462 = n461 ^ n459 ;
  assign n443 = x23 & ~x31 ;
  assign n450 = n176 & n443 ;
  assign n451 = n273 & n450 ;
  assign n448 = ~n260 & n443 ;
  assign n446 = n124 & n443 ;
  assign n444 = n170 & n443 ;
  assign n445 = n168 & n444 ;
  assign n447 = n446 ^ n445 ;
  assign n449 = n448 ^ n447 ;
  assign n452 = n451 ^ n449 ;
  assign n463 = n462 ^ n452 ;
  assign n467 = ~x30 & n463 ;
  assign n400 = x22 & n124 ;
  assign n403 = n402 ^ n400 ;
  assign n405 = n404 ^ n403 ;
  assign n408 = n407 ^ n405 ;
  assign n465 = n408 & n463 ;
  assign n391 = ~n124 & n236 ;
  assign n394 = n393 ^ n391 ;
  assign n396 = n395 ^ n394 ;
  assign n399 = n398 ^ n396 ;
  assign n464 = n399 & n463 ;
  assign n466 = n465 ^ n464 ;
  assign n468 = n467 ^ n466 ;
  assign n434 = x22 & ~x30 ;
  assign n440 = n176 & n434 ;
  assign n441 = n273 & n440 ;
  assign n438 = n434 & ~n437 ;
  assign n435 = n260 & n434 ;
  assign n439 = n438 ^ n435 ;
  assign n442 = n441 ^ n439 ;
  assign n469 = n468 ^ n442 ;
  assign n477 = n476 ^ n469 ;
  assign n478 = n390 & n477 ;
  assign n483 = n482 ^ n478 ;
  assign n484 = n349 & n483 ;
  assign n495 = n494 ^ n484 ;
  assign n409 = n408 ^ n399 ;
  assign n410 = n409 ^ x30 ;
  assign n420 = x23 & n124 ;
  assign n423 = n422 ^ n420 ;
  assign n425 = n424 ^ n423 ;
  assign n428 = n427 ^ n425 ;
  assign n411 = ~n124 & n256 ;
  assign n414 = n413 ^ n411 ;
  assign n416 = n415 ^ n414 ;
  assign n419 = n418 ^ n416 ;
  assign n429 = n428 ^ n419 ;
  assign n430 = n429 ^ x31 ;
  assign n431 = ~n410 & ~n430 ;
  assign n432 = n390 & n431 ;
  assign n433 = n349 & n432 ;
  assign n496 = n495 ^ n433 ;
  assign n877 = n285 & ~n496 ;
  assign n876 = x24 & n496 ;
  assign n878 = n877 ^ n876 ;
  assign n888 = n875 & ~n878 ;
  assign n879 = n878 ^ n875 ;
  assign n881 = n305 & ~n496 ;
  assign n880 = x25 & n496 ;
  assign n882 = n881 ^ n880 ;
  assign n884 = n699 & ~n872 ;
  assign n883 = n702 & n872 ;
  assign n885 = n884 ^ n883 ;
  assign n886 = ~n882 & n885 ;
  assign n887 = ~n879 & n886 ;
  assign n889 = n888 ^ n887 ;
  assign n1392 = n875 & n889 ;
  assign n892 = n326 & ~n496 ;
  assign n891 = x26 & n496 ;
  assign n893 = n892 ^ n891 ;
  assign n895 = n716 & ~n872 ;
  assign n894 = n707 & n872 ;
  assign n896 = n895 ^ n894 ;
  assign n906 = ~n893 & n896 ;
  assign n897 = n896 ^ n893 ;
  assign n899 = n729 & ~n872 ;
  assign n898 = n720 & n872 ;
  assign n900 = n899 ^ n898 ;
  assign n902 = n346 & ~n496 ;
  assign n901 = x27 & n496 ;
  assign n903 = n902 ^ n901 ;
  assign n904 = n900 & ~n903 ;
  assign n905 = ~n897 & n904 ;
  assign n907 = n906 ^ n905 ;
  assign n908 = n885 ^ n882 ;
  assign n909 = ~n879 & ~n908 ;
  assign n910 = n875 & n909 ;
  assign n911 = n907 & n910 ;
  assign n1393 = n1392 ^ n911 ;
  assign n913 = n903 ^ n900 ;
  assign n914 = ~n897 & ~n913 ;
  assign n915 = n909 & n914 ;
  assign n920 = n744 & ~n872 ;
  assign n919 = n735 & n872 ;
  assign n921 = n920 ^ n919 ;
  assign n917 = n368 & ~n496 ;
  assign n916 = x28 & n496 ;
  assign n918 = n917 ^ n916 ;
  assign n922 = n921 ^ n918 ;
  assign n927 = n757 & ~n872 ;
  assign n926 = n748 & n872 ;
  assign n928 = n927 ^ n926 ;
  assign n924 = n388 & ~n496 ;
  assign n923 = x29 & n496 ;
  assign n925 = n924 ^ n923 ;
  assign n929 = n928 ^ n925 ;
  assign n930 = ~n922 & ~n929 ;
  assign n935 = n768 & ~n872 ;
  assign n934 = n771 & n872 ;
  assign n936 = n935 ^ n934 ;
  assign n932 = n409 & ~n496 ;
  assign n931 = x30 & n496 ;
  assign n933 = n932 ^ n931 ;
  assign n937 = n936 ^ n933 ;
  assign n942 = n429 & ~n496 ;
  assign n941 = x31 & n496 ;
  assign n943 = n942 ^ n941 ;
  assign n939 = n781 & ~n872 ;
  assign n938 = n789 & n872 ;
  assign n940 = n939 ^ n938 ;
  assign n944 = n943 ^ n940 ;
  assign n945 = ~n937 & ~n944 ;
  assign n946 = n930 & n945 ;
  assign n947 = n915 & n946 ;
  assign n948 = n875 & ~n947 ;
  assign n1394 = n1393 ^ n948 ;
  assign n950 = n875 & n915 ;
  assign n958 = ~n918 & n921 ;
  assign n956 = ~n925 & n928 ;
  assign n957 = ~n922 & n956 ;
  assign n959 = n958 ^ n957 ;
  assign n953 = ~n933 & n936 ;
  assign n951 = n940 & ~n943 ;
  assign n952 = ~n937 & n951 ;
  assign n954 = n953 ^ n952 ;
  assign n955 = n930 & n954 ;
  assign n960 = n959 ^ n955 ;
  assign n961 = n950 & n960 ;
  assign n1395 = n1394 ^ n961 ;
  assign n1388 = n878 & ~n889 ;
  assign n964 = n878 & n909 ;
  assign n965 = n907 & n964 ;
  assign n1389 = n1388 ^ n965 ;
  assign n967 = n878 & ~n947 ;
  assign n1390 = n1389 ^ n967 ;
  assign n969 = n878 & n915 ;
  assign n970 = n960 & n969 ;
  assign n1391 = n1390 ^ n970 ;
  assign n1396 = n1395 ^ n1391 ;
  assign n1572 = ~n1396 & n1399 ;
  assign n1400 = n1399 ^ n1396 ;
  assign n1405 = n885 & n889 ;
  assign n975 = n885 & n909 ;
  assign n976 = n907 & n975 ;
  assign n1406 = n1405 ^ n976 ;
  assign n978 = n885 & ~n947 ;
  assign n1407 = n1406 ^ n978 ;
  assign n980 = n885 & n915 ;
  assign n981 = n960 & n980 ;
  assign n1408 = n1407 ^ n981 ;
  assign n1401 = n882 & ~n889 ;
  assign n984 = n882 & n909 ;
  assign n985 = n907 & n984 ;
  assign n1402 = n1401 ^ n985 ;
  assign n987 = n882 & ~n947 ;
  assign n1403 = n1402 ^ n987 ;
  assign n989 = n882 & n915 ;
  assign n990 = n960 & n989 ;
  assign n1404 = n1403 ^ n990 ;
  assign n1409 = n1408 ^ n1404 ;
  assign n1411 = n702 & ~n872 ;
  assign n1410 = n699 & n872 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1570 = ~n1409 & n1412 ;
  assign n1571 = ~n1400 & n1570 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1413 = n1412 ^ n1409 ;
  assign n1414 = ~n1400 & ~n1413 ;
  assign n1386 = n707 & ~n872 ;
  assign n1385 = n716 & n872 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1419 = n889 & n896 ;
  assign n1001 = n896 & n909 ;
  assign n1002 = n907 & n1001 ;
  assign n1420 = n1419 ^ n1002 ;
  assign n1004 = n896 & ~n947 ;
  assign n1421 = n1420 ^ n1004 ;
  assign n1006 = n896 & n915 ;
  assign n1007 = n960 & n1006 ;
  assign n1422 = n1421 ^ n1007 ;
  assign n1415 = ~n889 & n893 ;
  assign n1010 = n893 & n909 ;
  assign n1011 = n907 & n1010 ;
  assign n1416 = n1415 ^ n1011 ;
  assign n1013 = n893 & ~n947 ;
  assign n1417 = n1416 ^ n1013 ;
  assign n1015 = n893 & n915 ;
  assign n1016 = n960 & n1015 ;
  assign n1418 = n1417 ^ n1016 ;
  assign n1423 = n1422 ^ n1418 ;
  assign n1567 = n1387 & ~n1423 ;
  assign n1424 = n1423 ^ n1387 ;
  assign n1426 = n720 & ~n872 ;
  assign n1425 = n729 & n872 ;
  assign n1427 = n1426 ^ n1425 ;
  assign n1432 = n889 & n900 ;
  assign n1028 = n900 & n909 ;
  assign n1029 = n907 & n1028 ;
  assign n1433 = n1432 ^ n1029 ;
  assign n1031 = n900 & ~n947 ;
  assign n1434 = n1433 ^ n1031 ;
  assign n1033 = n900 & n915 ;
  assign n1034 = n960 & n1033 ;
  assign n1435 = n1434 ^ n1034 ;
  assign n1428 = ~n889 & n903 ;
  assign n1037 = n903 & n909 ;
  assign n1038 = n907 & n1037 ;
  assign n1429 = n1428 ^ n1038 ;
  assign n1040 = n903 & ~n947 ;
  assign n1430 = n1429 ^ n1040 ;
  assign n1042 = n903 & n915 ;
  assign n1043 = n960 & n1042 ;
  assign n1431 = n1430 ^ n1043 ;
  assign n1436 = n1435 ^ n1431 ;
  assign n1565 = n1427 & ~n1436 ;
  assign n1566 = ~n1424 & n1565 ;
  assign n1568 = n1567 ^ n1566 ;
  assign n1569 = n1414 & n1568 ;
  assign n1574 = n1573 ^ n1569 ;
  assign n1437 = n1436 ^ n1427 ;
  assign n1438 = ~n1424 & ~n1437 ;
  assign n1439 = n1414 & n1438 ;
  assign n1441 = n735 & ~n872 ;
  assign n1440 = n744 & n872 ;
  assign n1442 = n1441 ^ n1440 ;
  assign n1447 = n889 & n921 ;
  assign n1059 = n909 & n921 ;
  assign n1060 = n907 & n1059 ;
  assign n1448 = n1447 ^ n1060 ;
  assign n1062 = n921 & ~n947 ;
  assign n1449 = n1448 ^ n1062 ;
  assign n1064 = n915 & n921 ;
  assign n1065 = n960 & n1064 ;
  assign n1450 = n1449 ^ n1065 ;
  assign n1443 = ~n889 & n918 ;
  assign n1068 = n909 & n918 ;
  assign n1069 = n907 & n1068 ;
  assign n1444 = n1443 ^ n1069 ;
  assign n1071 = n918 & ~n947 ;
  assign n1445 = n1444 ^ n1071 ;
  assign n1073 = n915 & n918 ;
  assign n1074 = n960 & n1073 ;
  assign n1446 = n1445 ^ n1074 ;
  assign n1451 = n1450 ^ n1446 ;
  assign n1561 = n1442 & ~n1451 ;
  assign n1452 = n1451 ^ n1442 ;
  assign n1454 = n748 & ~n872 ;
  assign n1453 = n757 & n872 ;
  assign n1455 = n1454 ^ n1453 ;
  assign n1460 = n889 & n928 ;
  assign n1082 = n909 & n928 ;
  assign n1083 = n907 & n1082 ;
  assign n1461 = n1460 ^ n1083 ;
  assign n1085 = n928 & ~n947 ;
  assign n1462 = n1461 ^ n1085 ;
  assign n1087 = n915 & n928 ;
  assign n1088 = n960 & n1087 ;
  assign n1463 = n1462 ^ n1088 ;
  assign n1456 = ~n889 & n925 ;
  assign n1091 = n909 & n925 ;
  assign n1092 = n907 & n1091 ;
  assign n1457 = n1456 ^ n1092 ;
  assign n1094 = n925 & ~n947 ;
  assign n1458 = n1457 ^ n1094 ;
  assign n1096 = n915 & n925 ;
  assign n1097 = n960 & n1096 ;
  assign n1459 = n1458 ^ n1097 ;
  assign n1464 = n1463 ^ n1459 ;
  assign n1559 = n1455 & ~n1464 ;
  assign n1560 = ~n1452 & n1559 ;
  assign n1562 = n1561 ^ n1560 ;
  assign n1465 = n1464 ^ n1455 ;
  assign n1466 = ~n1452 & ~n1465 ;
  assign n1477 = n771 & ~n872 ;
  assign n1476 = n768 & n872 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1550 = ~n936 & n1478 ;
  assign n1554 = n915 & n1550 ;
  assign n1555 = n960 & n1554 ;
  assign n1496 = n907 & n909 ;
  assign n1497 = n1496 ^ n889 ;
  assign n1552 = ~n1497 & n1550 ;
  assign n1551 = n947 & n1550 ;
  assign n1553 = n1552 ^ n1551 ;
  assign n1556 = n1555 ^ n1553 ;
  assign n1490 = n789 & ~n872 ;
  assign n1489 = n781 & n872 ;
  assign n1491 = n1490 ^ n1489 ;
  assign n1515 = ~n943 & n1491 ;
  assign n1522 = n915 & n1515 ;
  assign n1523 = n960 & n1522 ;
  assign n1520 = ~n947 & n1515 ;
  assign n1518 = ~n889 & n1515 ;
  assign n1516 = n909 & n1515 ;
  assign n1517 = n907 & n1516 ;
  assign n1519 = n1518 ^ n1517 ;
  assign n1521 = n1520 ^ n1519 ;
  assign n1524 = n1523 ^ n1521 ;
  assign n1505 = ~n940 & n1491 ;
  assign n1512 = n915 & n1505 ;
  assign n1513 = n960 & n1512 ;
  assign n1510 = ~n947 & n1505 ;
  assign n1508 = n889 & n1505 ;
  assign n1506 = n909 & n1505 ;
  assign n1507 = n907 & n1506 ;
  assign n1509 = n1508 ^ n1507 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1514 = n1513 ^ n1511 ;
  assign n1525 = n1524 ^ n1514 ;
  assign n1547 = n1478 & n1525 ;
  assign n1542 = n915 & ~n936 ;
  assign n1543 = n960 & n1542 ;
  assign n1540 = ~n936 & ~n947 ;
  assign n1538 = n889 & ~n936 ;
  assign n1536 = n909 & ~n936 ;
  assign n1537 = n907 & n1536 ;
  assign n1539 = n1538 ^ n1537 ;
  assign n1541 = n1540 ^ n1539 ;
  assign n1544 = n1543 ^ n1541 ;
  assign n1545 = n1525 & n1544 ;
  assign n1532 = n915 & ~n933 ;
  assign n1533 = n960 & n1532 ;
  assign n1530 = ~n933 & ~n947 ;
  assign n1528 = ~n889 & ~n933 ;
  assign n1526 = n909 & ~n933 ;
  assign n1527 = n907 & n1526 ;
  assign n1529 = n1528 ^ n1527 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1534 = n1533 ^ n1531 ;
  assign n1535 = n1525 & n1534 ;
  assign n1546 = n1545 ^ n1535 ;
  assign n1548 = n1547 ^ n1546 ;
  assign n1498 = ~n933 & n1478 ;
  assign n1502 = n915 & n1498 ;
  assign n1503 = n960 & n1502 ;
  assign n1500 = ~n947 & n1498 ;
  assign n1499 = ~n1497 & n1498 ;
  assign n1501 = n1500 ^ n1499 ;
  assign n1504 = n1503 ^ n1501 ;
  assign n1549 = n1548 ^ n1504 ;
  assign n1557 = n1556 ^ n1549 ;
  assign n1558 = n1466 & n1557 ;
  assign n1563 = n1562 ^ n1558 ;
  assign n1564 = n1439 & n1563 ;
  assign n1575 = n1574 ^ n1564 ;
  assign n1471 = n889 & n936 ;
  assign n1106 = n909 & n936 ;
  assign n1107 = n907 & n1106 ;
  assign n1472 = n1471 ^ n1107 ;
  assign n1109 = n936 & ~n947 ;
  assign n1473 = n1472 ^ n1109 ;
  assign n1111 = n915 & n936 ;
  assign n1112 = n960 & n1111 ;
  assign n1474 = n1473 ^ n1112 ;
  assign n1467 = ~n889 & n933 ;
  assign n1115 = n909 & n933 ;
  assign n1116 = n907 & n1115 ;
  assign n1468 = n1467 ^ n1116 ;
  assign n1118 = n933 & ~n947 ;
  assign n1469 = n1468 ^ n1118 ;
  assign n1120 = n915 & n933 ;
  assign n1121 = n960 & n1120 ;
  assign n1470 = n1469 ^ n1121 ;
  assign n1475 = n1474 ^ n1470 ;
  assign n1479 = n1478 ^ n1475 ;
  assign n1484 = n889 & n940 ;
  assign n1132 = n909 & n940 ;
  assign n1133 = n907 & n1132 ;
  assign n1485 = n1484 ^ n1133 ;
  assign n1135 = n940 & ~n947 ;
  assign n1486 = n1485 ^ n1135 ;
  assign n1137 = n915 & n940 ;
  assign n1138 = n960 & n1137 ;
  assign n1487 = n1486 ^ n1138 ;
  assign n1480 = ~n889 & n943 ;
  assign n1141 = n909 & n943 ;
  assign n1142 = n907 & n1141 ;
  assign n1481 = n1480 ^ n1142 ;
  assign n1144 = n943 & ~n947 ;
  assign n1482 = n1481 ^ n1144 ;
  assign n1146 = n915 & n943 ;
  assign n1147 = n960 & n1146 ;
  assign n1483 = n1482 ^ n1147 ;
  assign n1488 = n1487 ^ n1483 ;
  assign n1492 = n1491 ^ n1488 ;
  assign n1493 = ~n1479 & ~n1492 ;
  assign n1494 = n1466 & n1493 ;
  assign n1495 = n1439 & n1494 ;
  assign n1576 = n1575 ^ n1495 ;
  assign n2040 = n1399 & ~n1576 ;
  assign n2039 = n1396 & n1576 ;
  assign n2041 = n2040 ^ n2039 ;
  assign n1607 = n1396 & ~n1576 ;
  assign n1606 = n1399 & n1576 ;
  assign n1608 = n1607 ^ n1606 ;
  assign n963 = n878 & n889 ;
  assign n966 = n965 ^ n963 ;
  assign n968 = n967 ^ n966 ;
  assign n971 = n970 ^ n968 ;
  assign n890 = n875 & ~n889 ;
  assign n912 = n911 ^ n890 ;
  assign n949 = n948 ^ n912 ;
  assign n962 = n961 ^ n949 ;
  assign n972 = n971 ^ n962 ;
  assign n498 = x24 & ~n496 ;
  assign n497 = n285 & n496 ;
  assign n499 = n498 ^ n497 ;
  assign n577 = ~x32 & n499 ;
  assign n500 = n499 ^ x32 ;
  assign n502 = x25 & ~n496 ;
  assign n501 = n305 & n496 ;
  assign n503 = n502 ^ n501 ;
  assign n575 = ~x33 & n503 ;
  assign n576 = ~n500 & n575 ;
  assign n578 = n577 ^ n576 ;
  assign n504 = n503 ^ x33 ;
  assign n505 = ~n500 & ~n504 ;
  assign n507 = x26 & ~n496 ;
  assign n506 = n326 & n496 ;
  assign n508 = n507 ^ n506 ;
  assign n572 = ~x34 & n508 ;
  assign n509 = n508 ^ x34 ;
  assign n568 = ~x35 & n346 ;
  assign n569 = n496 & n568 ;
  assign n566 = x27 & ~x35 ;
  assign n567 = ~n496 & n566 ;
  assign n570 = n569 ^ n567 ;
  assign n571 = ~n509 & n570 ;
  assign n573 = n572 ^ n571 ;
  assign n574 = n505 & n573 ;
  assign n579 = n578 ^ n574 ;
  assign n511 = x27 & ~n496 ;
  assign n510 = n346 & n496 ;
  assign n512 = n511 ^ n510 ;
  assign n513 = n512 ^ x35 ;
  assign n514 = ~n509 & ~n513 ;
  assign n515 = n505 & n514 ;
  assign n517 = x28 & ~n496 ;
  assign n516 = n368 & n496 ;
  assign n518 = n517 ^ n516 ;
  assign n562 = ~x36 & n518 ;
  assign n519 = n518 ^ x36 ;
  assign n558 = ~x37 & n388 ;
  assign n559 = n496 & n558 ;
  assign n556 = x29 & ~x37 ;
  assign n557 = ~n496 & n556 ;
  assign n560 = n559 ^ n557 ;
  assign n561 = ~n519 & n560 ;
  assign n563 = n562 ^ n561 ;
  assign n521 = x29 & ~n496 ;
  assign n520 = n388 & n496 ;
  assign n522 = n521 ^ n520 ;
  assign n523 = n522 ^ x37 ;
  assign n524 = ~n519 & ~n523 ;
  assign n552 = ~x38 & n409 ;
  assign n553 = n496 & n552 ;
  assign n541 = x31 & ~x39 ;
  assign n547 = ~x38 & n541 ;
  assign n548 = ~n496 & n547 ;
  assign n538 = ~x39 & n429 ;
  assign n545 = ~x38 & n538 ;
  assign n546 = n496 & n545 ;
  assign n549 = n548 ^ n546 ;
  assign n542 = x30 & n541 ;
  assign n543 = ~n496 & n542 ;
  assign n539 = n409 & n538 ;
  assign n540 = n496 & n539 ;
  assign n544 = n543 ^ n540 ;
  assign n550 = n549 ^ n544 ;
  assign n536 = x30 & ~x38 ;
  assign n537 = ~n496 & n536 ;
  assign n551 = n550 ^ n537 ;
  assign n554 = n553 ^ n551 ;
  assign n555 = n524 & n554 ;
  assign n564 = n563 ^ n555 ;
  assign n565 = n515 & n564 ;
  assign n580 = n579 ^ n565 ;
  assign n526 = x30 & ~n496 ;
  assign n525 = n409 & n496 ;
  assign n527 = n526 ^ n525 ;
  assign n528 = n527 ^ x38 ;
  assign n530 = x31 & ~n496 ;
  assign n529 = n429 & n496 ;
  assign n531 = n530 ^ n529 ;
  assign n532 = n531 ^ x39 ;
  assign n533 = ~n528 & ~n532 ;
  assign n534 = n524 & n533 ;
  assign n535 = n515 & n534 ;
  assign n581 = n580 ^ n535 ;
  assign n671 = n499 & ~n581 ;
  assign n670 = x32 & n581 ;
  assign n672 = n671 ^ n670 ;
  assign n998 = ~n672 & n972 ;
  assign n973 = n972 ^ n672 ;
  assign n983 = n882 & n889 ;
  assign n986 = n985 ^ n983 ;
  assign n988 = n987 ^ n986 ;
  assign n991 = n990 ^ n988 ;
  assign n974 = n885 & ~n889 ;
  assign n977 = n976 ^ n974 ;
  assign n979 = n978 ^ n977 ;
  assign n982 = n981 ^ n979 ;
  assign n992 = n991 ^ n982 ;
  assign n994 = n503 & ~n581 ;
  assign n993 = x33 & n581 ;
  assign n995 = n994 ^ n993 ;
  assign n996 = n992 & ~n995 ;
  assign n997 = ~n973 & n996 ;
  assign n999 = n998 ^ n997 ;
  assign n1613 = n972 & n999 ;
  assign n1009 = n889 & n893 ;
  assign n1012 = n1011 ^ n1009 ;
  assign n1014 = n1013 ^ n1012 ;
  assign n1017 = n1016 ^ n1014 ;
  assign n1000 = ~n889 & n896 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n1005 = n1004 ^ n1003 ;
  assign n1008 = n1007 ^ n1005 ;
  assign n1018 = n1017 ^ n1008 ;
  assign n1021 = n508 & ~n581 ;
  assign n1020 = x34 & n581 ;
  assign n1022 = n1021 ^ n1020 ;
  assign n1048 = n1018 & ~n1022 ;
  assign n1023 = n1022 ^ n1018 ;
  assign n1025 = n512 & ~n581 ;
  assign n1024 = x35 & n581 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1036 = n889 & n903 ;
  assign n1039 = n1038 ^ n1036 ;
  assign n1041 = n1040 ^ n1039 ;
  assign n1044 = n1043 ^ n1041 ;
  assign n1027 = ~n889 & n900 ;
  assign n1030 = n1029 ^ n1027 ;
  assign n1032 = n1031 ^ n1030 ;
  assign n1035 = n1034 ^ n1032 ;
  assign n1045 = n1044 ^ n1035 ;
  assign n1046 = ~n1026 & n1045 ;
  assign n1047 = ~n1023 & n1046 ;
  assign n1049 = n1048 ^ n1047 ;
  assign n1050 = n995 ^ n992 ;
  assign n1051 = ~n973 & ~n1050 ;
  assign n1210 = n972 & n1051 ;
  assign n1211 = n1049 & n1210 ;
  assign n1614 = n1613 ^ n1211 ;
  assign n1055 = n1045 ^ n1026 ;
  assign n1056 = ~n1023 & ~n1055 ;
  assign n1057 = n1051 & n1056 ;
  assign n1078 = n518 & ~n581 ;
  assign n1077 = x36 & n581 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1067 = n889 & n918 ;
  assign n1070 = n1069 ^ n1067 ;
  assign n1072 = n1071 ^ n1070 ;
  assign n1075 = n1074 ^ n1072 ;
  assign n1058 = ~n889 & n921 ;
  assign n1061 = n1060 ^ n1058 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1066 = n1065 ^ n1063 ;
  assign n1076 = n1075 ^ n1066 ;
  assign n1080 = n1079 ^ n1076 ;
  assign n1101 = n522 & ~n581 ;
  assign n1100 = x37 & n581 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1090 = n889 & n925 ;
  assign n1093 = n1092 ^ n1090 ;
  assign n1095 = n1094 ^ n1093 ;
  assign n1098 = n1097 ^ n1095 ;
  assign n1081 = ~n889 & n928 ;
  assign n1084 = n1083 ^ n1081 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1089 = n1088 ^ n1086 ;
  assign n1099 = n1098 ^ n1089 ;
  assign n1103 = n1102 ^ n1099 ;
  assign n1104 = ~n1080 & ~n1103 ;
  assign n1125 = n527 & ~n581 ;
  assign n1124 = x38 & n581 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1114 = n889 & n933 ;
  assign n1117 = n1116 ^ n1114 ;
  assign n1119 = n1118 ^ n1117 ;
  assign n1122 = n1121 ^ n1119 ;
  assign n1105 = ~n889 & n936 ;
  assign n1108 = n1107 ^ n1105 ;
  assign n1110 = n1109 ^ n1108 ;
  assign n1113 = n1112 ^ n1110 ;
  assign n1123 = n1122 ^ n1113 ;
  assign n1127 = n1126 ^ n1123 ;
  assign n1140 = n889 & n943 ;
  assign n1143 = n1142 ^ n1140 ;
  assign n1145 = n1144 ^ n1143 ;
  assign n1148 = n1147 ^ n1145 ;
  assign n1131 = ~n889 & n940 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1139 = n1138 ^ n1136 ;
  assign n1149 = n1148 ^ n1139 ;
  assign n1129 = n531 & ~n581 ;
  assign n1128 = x39 & n581 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1150 = n1149 ^ n1130 ;
  assign n1151 = ~n1127 & ~n1150 ;
  assign n1152 = n1104 & n1151 ;
  assign n1153 = n1057 & n1152 ;
  assign n1213 = n972 & ~n1153 ;
  assign n1615 = n1614 ^ n1213 ;
  assign n1163 = n1076 & ~n1079 ;
  assign n1161 = n1099 & ~n1102 ;
  assign n1162 = ~n1080 & n1161 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n1158 = n1123 & ~n1126 ;
  assign n1156 = ~n1130 & n1149 ;
  assign n1157 = ~n1127 & n1156 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1160 = n1104 & n1159 ;
  assign n1165 = n1164 ^ n1160 ;
  assign n1215 = n972 & n1057 ;
  assign n1216 = n1165 & n1215 ;
  assign n1616 = n1615 ^ n1216 ;
  assign n1609 = n672 & ~n999 ;
  assign n1219 = n672 & n1051 ;
  assign n1220 = n1049 & n1219 ;
  assign n1610 = n1609 ^ n1220 ;
  assign n1222 = n672 & ~n1153 ;
  assign n1611 = n1610 ^ n1222 ;
  assign n1224 = n672 & n1057 ;
  assign n1225 = n1165 & n1224 ;
  assign n1612 = n1611 ^ n1225 ;
  assign n1617 = n1616 ^ n1612 ;
  assign n1637 = n1608 & ~n1617 ;
  assign n1618 = n1617 ^ n1608 ;
  assign n1623 = n992 & n999 ;
  assign n1233 = n992 & n1051 ;
  assign n1234 = n1049 & n1233 ;
  assign n1624 = n1623 ^ n1234 ;
  assign n1236 = n992 & ~n1153 ;
  assign n1625 = n1624 ^ n1236 ;
  assign n1238 = n992 & n1057 ;
  assign n1239 = n1165 & n1238 ;
  assign n1626 = n1625 ^ n1239 ;
  assign n1619 = n995 & ~n999 ;
  assign n1242 = n995 & n1051 ;
  assign n1243 = n1049 & n1242 ;
  assign n1620 = n1619 ^ n1243 ;
  assign n1245 = n995 & ~n1153 ;
  assign n1621 = n1620 ^ n1245 ;
  assign n1247 = n995 & n1057 ;
  assign n1248 = n1165 & n1247 ;
  assign n1622 = n1621 ^ n1248 ;
  assign n1627 = n1626 ^ n1622 ;
  assign n1629 = n1409 & ~n1576 ;
  assign n1628 = n1412 & n1576 ;
  assign n1630 = n1629 ^ n1628 ;
  assign n1635 = ~n1627 & n1630 ;
  assign n1636 = ~n1618 & n1635 ;
  assign n1638 = n1637 ^ n1636 ;
  assign n2046 = n1608 & n1638 ;
  assign n1578 = n1423 & ~n1576 ;
  assign n1577 = n1387 & n1576 ;
  assign n1579 = n1578 ^ n1577 ;
  assign n1584 = n999 & n1018 ;
  assign n1052 = n1018 & n1051 ;
  assign n1053 = n1049 & n1052 ;
  assign n1585 = n1584 ^ n1053 ;
  assign n1154 = n1018 & ~n1153 ;
  assign n1586 = n1585 ^ n1154 ;
  assign n1166 = n1018 & n1057 ;
  assign n1167 = n1165 & n1166 ;
  assign n1587 = n1586 ^ n1167 ;
  assign n1580 = ~n999 & n1022 ;
  assign n1170 = n1022 & n1051 ;
  assign n1171 = n1049 & n1170 ;
  assign n1581 = n1580 ^ n1171 ;
  assign n1173 = n1022 & ~n1153 ;
  assign n1582 = n1581 ^ n1173 ;
  assign n1175 = n1022 & n1057 ;
  assign n1176 = n1165 & n1175 ;
  assign n1583 = n1582 ^ n1176 ;
  assign n1588 = n1587 ^ n1583 ;
  assign n1604 = n1579 & ~n1588 ;
  assign n1589 = n1588 ^ n1579 ;
  assign n1591 = n1436 & ~n1576 ;
  assign n1590 = n1427 & n1576 ;
  assign n1592 = n1591 ^ n1590 ;
  assign n1597 = n999 & n1045 ;
  assign n1184 = n1045 & n1051 ;
  assign n1185 = n1049 & n1184 ;
  assign n1598 = n1597 ^ n1185 ;
  assign n1187 = n1045 & ~n1153 ;
  assign n1599 = n1598 ^ n1187 ;
  assign n1189 = n1045 & n1057 ;
  assign n1190 = n1165 & n1189 ;
  assign n1600 = n1599 ^ n1190 ;
  assign n1593 = ~n999 & n1026 ;
  assign n1193 = n1026 & n1051 ;
  assign n1194 = n1049 & n1193 ;
  assign n1594 = n1593 ^ n1194 ;
  assign n1196 = n1026 & ~n1153 ;
  assign n1595 = n1594 ^ n1196 ;
  assign n1198 = n1026 & n1057 ;
  assign n1199 = n1165 & n1198 ;
  assign n1596 = n1595 ^ n1199 ;
  assign n1601 = n1600 ^ n1596 ;
  assign n1602 = n1592 & ~n1601 ;
  assign n1603 = ~n1589 & n1602 ;
  assign n1605 = n1604 ^ n1603 ;
  assign n1631 = n1630 ^ n1627 ;
  assign n1632 = ~n1618 & ~n1631 ;
  assign n1633 = n1608 & n1632 ;
  assign n1634 = n1605 & n1633 ;
  assign n2047 = n2046 ^ n1634 ;
  assign n1641 = n1601 ^ n1592 ;
  assign n1642 = ~n1589 & ~n1641 ;
  assign n1643 = n1632 & n1642 ;
  assign n1654 = n1451 & ~n1576 ;
  assign n1653 = n1442 & n1576 ;
  assign n1655 = n1654 ^ n1653 ;
  assign n1648 = n999 & n1076 ;
  assign n1265 = n1051 & n1076 ;
  assign n1266 = n1049 & n1265 ;
  assign n1649 = n1648 ^ n1266 ;
  assign n1268 = n1076 & ~n1153 ;
  assign n1650 = n1649 ^ n1268 ;
  assign n1270 = n1057 & n1076 ;
  assign n1271 = n1165 & n1270 ;
  assign n1651 = n1650 ^ n1271 ;
  assign n1644 = ~n999 & n1079 ;
  assign n1274 = n1051 & n1079 ;
  assign n1275 = n1049 & n1274 ;
  assign n1645 = n1644 ^ n1275 ;
  assign n1277 = n1079 & ~n1153 ;
  assign n1646 = n1645 ^ n1277 ;
  assign n1279 = n1057 & n1079 ;
  assign n1280 = n1165 & n1279 ;
  assign n1647 = n1646 ^ n1280 ;
  assign n1652 = n1651 ^ n1647 ;
  assign n1656 = n1655 ^ n1652 ;
  assign n1667 = n1464 & ~n1576 ;
  assign n1666 = n1455 & n1576 ;
  assign n1668 = n1667 ^ n1666 ;
  assign n1661 = n999 & n1099 ;
  assign n1288 = n1051 & n1099 ;
  assign n1289 = n1049 & n1288 ;
  assign n1662 = n1661 ^ n1289 ;
  assign n1291 = n1099 & ~n1153 ;
  assign n1663 = n1662 ^ n1291 ;
  assign n1293 = n1057 & n1099 ;
  assign n1294 = n1165 & n1293 ;
  assign n1664 = n1663 ^ n1294 ;
  assign n1657 = ~n999 & n1102 ;
  assign n1297 = n1051 & n1102 ;
  assign n1298 = n1049 & n1297 ;
  assign n1658 = n1657 ^ n1298 ;
  assign n1300 = n1102 & ~n1153 ;
  assign n1659 = n1658 ^ n1300 ;
  assign n1302 = n1057 & n1102 ;
  assign n1303 = n1165 & n1302 ;
  assign n1660 = n1659 ^ n1303 ;
  assign n1665 = n1664 ^ n1660 ;
  assign n1669 = n1668 ^ n1665 ;
  assign n1670 = ~n1656 & ~n1669 ;
  assign n1681 = n1475 & ~n1576 ;
  assign n1680 = n1478 & n1576 ;
  assign n1682 = n1681 ^ n1680 ;
  assign n1675 = n999 & n1123 ;
  assign n1312 = n1051 & n1123 ;
  assign n1313 = n1049 & n1312 ;
  assign n1676 = n1675 ^ n1313 ;
  assign n1315 = n1123 & ~n1153 ;
  assign n1677 = n1676 ^ n1315 ;
  assign n1317 = n1057 & n1123 ;
  assign n1318 = n1165 & n1317 ;
  assign n1678 = n1677 ^ n1318 ;
  assign n1671 = ~n999 & n1126 ;
  assign n1321 = n1051 & n1126 ;
  assign n1322 = n1049 & n1321 ;
  assign n1672 = n1671 ^ n1322 ;
  assign n1324 = n1126 & ~n1153 ;
  assign n1673 = n1672 ^ n1324 ;
  assign n1326 = n1057 & n1126 ;
  assign n1327 = n1165 & n1326 ;
  assign n1674 = n1673 ^ n1327 ;
  assign n1679 = n1678 ^ n1674 ;
  assign n1683 = n1682 ^ n1679 ;
  assign n1691 = n999 & n1149 ;
  assign n1335 = n1051 & n1149 ;
  assign n1336 = n1049 & n1335 ;
  assign n1692 = n1691 ^ n1336 ;
  assign n1338 = n1149 & ~n1153 ;
  assign n1693 = n1692 ^ n1338 ;
  assign n1340 = n1057 & n1149 ;
  assign n1341 = n1165 & n1340 ;
  assign n1694 = n1693 ^ n1341 ;
  assign n1687 = ~n999 & n1130 ;
  assign n1344 = n1051 & n1130 ;
  assign n1345 = n1049 & n1344 ;
  assign n1688 = n1687 ^ n1345 ;
  assign n1347 = n1130 & ~n1153 ;
  assign n1689 = n1688 ^ n1347 ;
  assign n1349 = n1057 & n1130 ;
  assign n1350 = n1165 & n1349 ;
  assign n1690 = n1689 ^ n1350 ;
  assign n1695 = n1694 ^ n1690 ;
  assign n1685 = n1488 & ~n1576 ;
  assign n1684 = n1491 & n1576 ;
  assign n1686 = n1685 ^ n1684 ;
  assign n1696 = n1695 ^ n1686 ;
  assign n1697 = ~n1683 & ~n1696 ;
  assign n1698 = n1670 & n1697 ;
  assign n1699 = n1643 & n1698 ;
  assign n1700 = n1608 & ~n1699 ;
  assign n2048 = n2047 ^ n1700 ;
  assign n1702 = n1608 & n1643 ;
  assign n1710 = ~n1652 & n1655 ;
  assign n1708 = ~n1665 & n1668 ;
  assign n1709 = ~n1656 & n1708 ;
  assign n1711 = n1710 ^ n1709 ;
  assign n1705 = ~n1679 & n1682 ;
  assign n1703 = n1686 & ~n1695 ;
  assign n1704 = ~n1683 & n1703 ;
  assign n1706 = n1705 ^ n1704 ;
  assign n1707 = n1670 & n1706 ;
  assign n1712 = n1711 ^ n1707 ;
  assign n1713 = n1702 & n1712 ;
  assign n2049 = n2048 ^ n1713 ;
  assign n2042 = n1617 & ~n1638 ;
  assign n1715 = n1617 & n1632 ;
  assign n1716 = n1605 & n1715 ;
  assign n2043 = n2042 ^ n1716 ;
  assign n1719 = n1617 & ~n1699 ;
  assign n2044 = n2043 ^ n1719 ;
  assign n1721 = n1617 & n1643 ;
  assign n1722 = n1712 & n1721 ;
  assign n2045 = n2044 ^ n1722 ;
  assign n2050 = n2049 ^ n2045 ;
  assign n2226 = n2041 & ~n2050 ;
  assign n2051 = n2050 ^ n2041 ;
  assign n2056 = n1630 & n1638 ;
  assign n1726 = n1630 & n1632 ;
  assign n1727 = n1605 & n1726 ;
  assign n2057 = n2056 ^ n1727 ;
  assign n1730 = n1630 & ~n1699 ;
  assign n2058 = n2057 ^ n1730 ;
  assign n1732 = n1630 & n1643 ;
  assign n1733 = n1712 & n1732 ;
  assign n2059 = n2058 ^ n1733 ;
  assign n2052 = n1627 & ~n1638 ;
  assign n1735 = n1627 & n1632 ;
  assign n1736 = n1605 & n1735 ;
  assign n2053 = n2052 ^ n1736 ;
  assign n1739 = n1627 & ~n1699 ;
  assign n2054 = n2053 ^ n1739 ;
  assign n1741 = n1627 & n1643 ;
  assign n1742 = n1712 & n1741 ;
  assign n2055 = n2054 ^ n1742 ;
  assign n2060 = n2059 ^ n2055 ;
  assign n2062 = n1412 & ~n1576 ;
  assign n2061 = n1409 & n1576 ;
  assign n2063 = n2062 ^ n2061 ;
  assign n2224 = ~n2060 & n2063 ;
  assign n2225 = ~n2051 & n2224 ;
  assign n2227 = n2226 ^ n2225 ;
  assign n2064 = n2063 ^ n2060 ;
  assign n2065 = ~n2051 & ~n2064 ;
  assign n2067 = n1387 & ~n1576 ;
  assign n2066 = n1423 & n1576 ;
  assign n2068 = n2067 ^ n2066 ;
  assign n2073 = n1579 & n1638 ;
  assign n1766 = n1579 & n1632 ;
  assign n1767 = n1605 & n1766 ;
  assign n2074 = n2073 ^ n1767 ;
  assign n1770 = n1579 & ~n1699 ;
  assign n2075 = n2074 ^ n1770 ;
  assign n1772 = n1579 & n1643 ;
  assign n1773 = n1712 & n1772 ;
  assign n2076 = n2075 ^ n1773 ;
  assign n2069 = n1588 & ~n1638 ;
  assign n1775 = n1588 & n1632 ;
  assign n1776 = n1605 & n1775 ;
  assign n2070 = n2069 ^ n1776 ;
  assign n1779 = n1588 & ~n1699 ;
  assign n2071 = n2070 ^ n1779 ;
  assign n1781 = n1588 & n1643 ;
  assign n1782 = n1712 & n1781 ;
  assign n2072 = n2071 ^ n1782 ;
  assign n2077 = n2076 ^ n2072 ;
  assign n2221 = n2068 & ~n2077 ;
  assign n2078 = n2077 ^ n2068 ;
  assign n2080 = n1427 & ~n1576 ;
  assign n2079 = n1436 & n1576 ;
  assign n2081 = n2080 ^ n2079 ;
  assign n2086 = n1592 & n1638 ;
  assign n1824 = n1592 & n1632 ;
  assign n1825 = n1605 & n1824 ;
  assign n2087 = n2086 ^ n1825 ;
  assign n1828 = n1592 & ~n1699 ;
  assign n2088 = n2087 ^ n1828 ;
  assign n1830 = n1592 & n1643 ;
  assign n1831 = n1712 & n1830 ;
  assign n2089 = n2088 ^ n1831 ;
  assign n2082 = n1601 & ~n1638 ;
  assign n1833 = n1601 & n1632 ;
  assign n1834 = n1605 & n1833 ;
  assign n2083 = n2082 ^ n1834 ;
  assign n1837 = n1601 & ~n1699 ;
  assign n2084 = n2083 ^ n1837 ;
  assign n1839 = n1601 & n1643 ;
  assign n1840 = n1712 & n1839 ;
  assign n2085 = n2084 ^ n1840 ;
  assign n2090 = n2089 ^ n2085 ;
  assign n2219 = n2081 & ~n2090 ;
  assign n2220 = ~n2078 & n2219 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2223 = n2065 & n2222 ;
  assign n2228 = n2227 ^ n2223 ;
  assign n2091 = n2090 ^ n2081 ;
  assign n2092 = ~n2078 & ~n2091 ;
  assign n2093 = n2065 & n2092 ;
  assign n2095 = n1442 & ~n1576 ;
  assign n2094 = n1451 & n1576 ;
  assign n2096 = n2095 ^ n2094 ;
  assign n2101 = n1638 & n1655 ;
  assign n1857 = n1632 & n1655 ;
  assign n1858 = n1605 & n1857 ;
  assign n2102 = n2101 ^ n1858 ;
  assign n1861 = n1655 & ~n1699 ;
  assign n2103 = n2102 ^ n1861 ;
  assign n1863 = n1643 & n1655 ;
  assign n1864 = n1712 & n1863 ;
  assign n2104 = n2103 ^ n1864 ;
  assign n2097 = ~n1638 & n1652 ;
  assign n1866 = n1632 & n1652 ;
  assign n1867 = n1605 & n1866 ;
  assign n2098 = n2097 ^ n1867 ;
  assign n1870 = n1652 & ~n1699 ;
  assign n2099 = n2098 ^ n1870 ;
  assign n1872 = n1643 & n1652 ;
  assign n1873 = n1712 & n1872 ;
  assign n2100 = n2099 ^ n1873 ;
  assign n2105 = n2104 ^ n2100 ;
  assign n2215 = n2096 & ~n2105 ;
  assign n2106 = n2105 ^ n2096 ;
  assign n2108 = n1455 & ~n1576 ;
  assign n2107 = n1464 & n1576 ;
  assign n2109 = n2108 ^ n2107 ;
  assign n2114 = n1638 & n1668 ;
  assign n1896 = n1632 & n1668 ;
  assign n1897 = n1605 & n1896 ;
  assign n2115 = n2114 ^ n1897 ;
  assign n1900 = n1668 & ~n1699 ;
  assign n2116 = n2115 ^ n1900 ;
  assign n1902 = n1643 & n1668 ;
  assign n1903 = n1712 & n1902 ;
  assign n2117 = n2116 ^ n1903 ;
  assign n2110 = ~n1638 & n1665 ;
  assign n1905 = n1632 & n1665 ;
  assign n1906 = n1605 & n1905 ;
  assign n2111 = n2110 ^ n1906 ;
  assign n1909 = n1665 & ~n1699 ;
  assign n2112 = n2111 ^ n1909 ;
  assign n1911 = n1643 & n1665 ;
  assign n1912 = n1712 & n1911 ;
  assign n2113 = n2112 ^ n1912 ;
  assign n2118 = n2117 ^ n2113 ;
  assign n2213 = n2109 & ~n2118 ;
  assign n2214 = ~n2106 & n2213 ;
  assign n2216 = n2215 ^ n2214 ;
  assign n2119 = n2118 ^ n2109 ;
  assign n2120 = ~n2106 & ~n2119 ;
  assign n2131 = n1478 & ~n1576 ;
  assign n2130 = n1475 & n1576 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2204 = ~n1682 & n2132 ;
  assign n2208 = n1643 & n2204 ;
  assign n2209 = n1712 & n2208 ;
  assign n2150 = n1605 & n1632 ;
  assign n2151 = n2150 ^ n1638 ;
  assign n2206 = ~n2151 & n2204 ;
  assign n2205 = n1699 & n2204 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2210 = n2209 ^ n2207 ;
  assign n2144 = n1491 & ~n1576 ;
  assign n2143 = n1488 & n1576 ;
  assign n2145 = n2144 ^ n2143 ;
  assign n2169 = ~n1695 & n2145 ;
  assign n2176 = n1643 & n2169 ;
  assign n2177 = n1712 & n2176 ;
  assign n2174 = ~n1699 & n2169 ;
  assign n2172 = ~n1638 & n2169 ;
  assign n2170 = n1632 & n2169 ;
  assign n2171 = n1605 & n2170 ;
  assign n2173 = n2172 ^ n2171 ;
  assign n2175 = n2174 ^ n2173 ;
  assign n2178 = n2177 ^ n2175 ;
  assign n2159 = ~n1686 & n2145 ;
  assign n2166 = n1643 & n2159 ;
  assign n2167 = n1712 & n2166 ;
  assign n2164 = ~n1699 & n2159 ;
  assign n2162 = n1638 & n2159 ;
  assign n2160 = n1632 & n2159 ;
  assign n2161 = n1605 & n2160 ;
  assign n2163 = n2162 ^ n2161 ;
  assign n2165 = n2164 ^ n2163 ;
  assign n2168 = n2167 ^ n2165 ;
  assign n2179 = n2178 ^ n2168 ;
  assign n2201 = n2132 & n2179 ;
  assign n2196 = n1643 & ~n1682 ;
  assign n2197 = n1712 & n2196 ;
  assign n2194 = ~n1682 & ~n1699 ;
  assign n2192 = n1638 & ~n1682 ;
  assign n2190 = n1632 & ~n1682 ;
  assign n2191 = n1605 & n2190 ;
  assign n2193 = n2192 ^ n2191 ;
  assign n2195 = n2194 ^ n2193 ;
  assign n2198 = n2197 ^ n2195 ;
  assign n2199 = n2179 & n2198 ;
  assign n2186 = n1643 & ~n1679 ;
  assign n2187 = n1712 & n2186 ;
  assign n2184 = ~n1679 & ~n1699 ;
  assign n2182 = ~n1638 & ~n1679 ;
  assign n2180 = n1632 & ~n1679 ;
  assign n2181 = n1605 & n2180 ;
  assign n2183 = n2182 ^ n2181 ;
  assign n2185 = n2184 ^ n2183 ;
  assign n2188 = n2187 ^ n2185 ;
  assign n2189 = n2179 & n2188 ;
  assign n2200 = n2199 ^ n2189 ;
  assign n2202 = n2201 ^ n2200 ;
  assign n2152 = ~n1679 & n2132 ;
  assign n2156 = n1643 & n2152 ;
  assign n2157 = n1712 & n2156 ;
  assign n2154 = ~n1699 & n2152 ;
  assign n2153 = ~n2151 & n2152 ;
  assign n2155 = n2154 ^ n2153 ;
  assign n2158 = n2157 ^ n2155 ;
  assign n2203 = n2202 ^ n2158 ;
  assign n2211 = n2210 ^ n2203 ;
  assign n2212 = n2120 & n2211 ;
  assign n2217 = n2216 ^ n2212 ;
  assign n2218 = n2093 & n2217 ;
  assign n2229 = n2228 ^ n2218 ;
  assign n2125 = n1638 & n1682 ;
  assign n1936 = n1632 & n1682 ;
  assign n1937 = n1605 & n1936 ;
  assign n2126 = n2125 ^ n1937 ;
  assign n1940 = n1682 & ~n1699 ;
  assign n2127 = n2126 ^ n1940 ;
  assign n1942 = n1643 & n1682 ;
  assign n1943 = n1712 & n1942 ;
  assign n2128 = n2127 ^ n1943 ;
  assign n2121 = ~n1638 & n1679 ;
  assign n1945 = n1632 & n1679 ;
  assign n1946 = n1605 & n1945 ;
  assign n2122 = n2121 ^ n1946 ;
  assign n1949 = n1679 & ~n1699 ;
  assign n2123 = n2122 ^ n1949 ;
  assign n1951 = n1643 & n1679 ;
  assign n1952 = n1712 & n1951 ;
  assign n2124 = n2123 ^ n1952 ;
  assign n2129 = n2128 ^ n2124 ;
  assign n2133 = n2132 ^ n2129 ;
  assign n2138 = n1638 & n1686 ;
  assign n1975 = n1632 & n1686 ;
  assign n1976 = n1605 & n1975 ;
  assign n2139 = n2138 ^ n1976 ;
  assign n1979 = n1686 & ~n1699 ;
  assign n2140 = n2139 ^ n1979 ;
  assign n1981 = n1643 & n1686 ;
  assign n1982 = n1712 & n1981 ;
  assign n2141 = n2140 ^ n1982 ;
  assign n2134 = ~n1638 & n1695 ;
  assign n1984 = n1632 & n1695 ;
  assign n1985 = n1605 & n1984 ;
  assign n2135 = n2134 ^ n1985 ;
  assign n1988 = n1695 & ~n1699 ;
  assign n2136 = n2135 ^ n1988 ;
  assign n1990 = n1643 & n1695 ;
  assign n1991 = n1712 & n1990 ;
  assign n2137 = n2136 ^ n1991 ;
  assign n2142 = n2141 ^ n2137 ;
  assign n2146 = n2145 ^ n2142 ;
  assign n2147 = ~n2133 & ~n2146 ;
  assign n2148 = n2120 & n2147 ;
  assign n2149 = n2093 & n2148 ;
  assign n2230 = n2229 ^ n2149 ;
  assign n2401 = n2041 & ~n2230 ;
  assign n2400 = n2050 & n2230 ;
  assign n2402 = n2401 ^ n2400 ;
  assign n2301 = n2105 & ~n2230 ;
  assign n2300 = n2096 & n2230 ;
  assign n2302 = n2301 ^ n2300 ;
  assign n1868 = n1638 & n1652 ;
  assign n1869 = n1868 ^ n1867 ;
  assign n1871 = n1870 ^ n1869 ;
  assign n1874 = n1873 ^ n1871 ;
  assign n1859 = ~n1638 & n1655 ;
  assign n1860 = n1859 ^ n1858 ;
  assign n1862 = n1861 ^ n1860 ;
  assign n1865 = n1864 ^ n1862 ;
  assign n1875 = n1874 ^ n1865 ;
  assign n1273 = n999 & n1079 ;
  assign n1276 = n1275 ^ n1273 ;
  assign n1278 = n1277 ^ n1276 ;
  assign n1281 = n1280 ^ n1278 ;
  assign n1264 = ~n999 & n1076 ;
  assign n1267 = n1266 ^ n1264 ;
  assign n1269 = n1268 ^ n1267 ;
  assign n1272 = n1271 ^ n1269 ;
  assign n1282 = n1281 ^ n1272 ;
  assign n602 = x36 & ~n581 ;
  assign n601 = n518 & n581 ;
  assign n603 = n602 ^ n601 ;
  assign n583 = x32 & ~n581 ;
  assign n582 = n499 & n581 ;
  assign n584 = n583 ^ n582 ;
  assign n662 = ~x40 & n584 ;
  assign n585 = n584 ^ x40 ;
  assign n587 = x33 & ~n581 ;
  assign n586 = n503 & n581 ;
  assign n588 = n587 ^ n586 ;
  assign n660 = ~x41 & n588 ;
  assign n661 = ~n585 & n660 ;
  assign n663 = n662 ^ n661 ;
  assign n589 = n588 ^ x41 ;
  assign n590 = ~n585 & ~n589 ;
  assign n592 = x34 & ~n581 ;
  assign n591 = n508 & n581 ;
  assign n593 = n592 ^ n591 ;
  assign n657 = ~x42 & n593 ;
  assign n594 = n593 ^ x42 ;
  assign n653 = ~x43 & n512 ;
  assign n654 = n581 & n653 ;
  assign n651 = x35 & ~x43 ;
  assign n652 = ~n581 & n651 ;
  assign n655 = n654 ^ n652 ;
  assign n656 = ~n594 & n655 ;
  assign n658 = n657 ^ n656 ;
  assign n659 = n590 & n658 ;
  assign n664 = n663 ^ n659 ;
  assign n596 = x35 & ~n581 ;
  assign n595 = n512 & n581 ;
  assign n597 = n596 ^ n595 ;
  assign n598 = n597 ^ x43 ;
  assign n599 = ~n594 & ~n598 ;
  assign n600 = n590 & n599 ;
  assign n647 = ~x44 & n603 ;
  assign n604 = n603 ^ x44 ;
  assign n643 = ~x45 & n522 ;
  assign n644 = n581 & n643 ;
  assign n641 = x37 & ~x45 ;
  assign n642 = ~n581 & n641 ;
  assign n645 = n644 ^ n642 ;
  assign n646 = ~n604 & n645 ;
  assign n648 = n647 ^ n646 ;
  assign n606 = x37 & ~n581 ;
  assign n605 = n522 & n581 ;
  assign n607 = n606 ^ n605 ;
  assign n608 = n607 ^ x45 ;
  assign n609 = ~n604 & ~n608 ;
  assign n637 = ~x46 & n527 ;
  assign n638 = n581 & n637 ;
  assign n626 = x39 & ~x47 ;
  assign n632 = ~x46 & n626 ;
  assign n633 = ~n581 & n632 ;
  assign n623 = ~x47 & n531 ;
  assign n630 = ~x46 & n623 ;
  assign n631 = n581 & n630 ;
  assign n634 = n633 ^ n631 ;
  assign n627 = x38 & n626 ;
  assign n628 = ~n581 & n627 ;
  assign n624 = n527 & n623 ;
  assign n625 = n581 & n624 ;
  assign n629 = n628 ^ n625 ;
  assign n635 = n634 ^ n629 ;
  assign n621 = x38 & ~x46 ;
  assign n622 = ~n581 & n621 ;
  assign n636 = n635 ^ n622 ;
  assign n639 = n638 ^ n636 ;
  assign n640 = n609 & n639 ;
  assign n649 = n648 ^ n640 ;
  assign n650 = n600 & n649 ;
  assign n665 = n664 ^ n650 ;
  assign n611 = x38 & ~n581 ;
  assign n610 = n527 & n581 ;
  assign n612 = n611 ^ n610 ;
  assign n613 = n612 ^ x46 ;
  assign n615 = x39 & ~n581 ;
  assign n614 = n531 & n581 ;
  assign n616 = n615 ^ n614 ;
  assign n617 = n616 ^ x47 ;
  assign n618 = ~n613 & ~n617 ;
  assign n619 = n609 & n618 ;
  assign n620 = n600 & n619 ;
  assign n666 = n665 ^ n620 ;
  assign n1284 = n603 & ~n666 ;
  assign n1283 = x44 & n666 ;
  assign n1285 = n1284 ^ n1283 ;
  assign n1369 = n1282 & ~n1285 ;
  assign n1286 = n1285 ^ n1282 ;
  assign n1296 = n999 & n1102 ;
  assign n1299 = n1298 ^ n1296 ;
  assign n1301 = n1300 ^ n1299 ;
  assign n1304 = n1303 ^ n1301 ;
  assign n1287 = ~n999 & n1099 ;
  assign n1290 = n1289 ^ n1287 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1295 = n1294 ^ n1292 ;
  assign n1305 = n1304 ^ n1295 ;
  assign n1307 = n607 & ~n666 ;
  assign n1306 = x45 & n666 ;
  assign n1308 = n1307 ^ n1306 ;
  assign n1367 = n1305 & ~n1308 ;
  assign n1368 = ~n1286 & n1367 ;
  assign n1370 = n1369 ^ n1368 ;
  assign n1309 = n1308 ^ n1305 ;
  assign n1310 = ~n1286 & ~n1309 ;
  assign n1320 = n999 & n1126 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1328 = n1327 ^ n1325 ;
  assign n1311 = ~n999 & n1123 ;
  assign n1314 = n1313 ^ n1311 ;
  assign n1316 = n1315 ^ n1314 ;
  assign n1319 = n1318 ^ n1316 ;
  assign n1329 = n1328 ^ n1319 ;
  assign n1331 = n612 & ~n666 ;
  assign n1330 = x46 & n666 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1364 = n1329 & ~n1332 ;
  assign n1333 = n1332 ^ n1329 ;
  assign n1343 = n999 & n1130 ;
  assign n1346 = n1345 ^ n1343 ;
  assign n1348 = n1347 ^ n1346 ;
  assign n1351 = n1350 ^ n1348 ;
  assign n1334 = ~n999 & n1149 ;
  assign n1337 = n1336 ^ n1334 ;
  assign n1339 = n1338 ^ n1337 ;
  assign n1342 = n1341 ^ n1339 ;
  assign n1352 = n1351 ^ n1342 ;
  assign n1354 = n616 & ~n666 ;
  assign n1353 = x47 & n666 ;
  assign n1355 = n1354 ^ n1353 ;
  assign n1362 = n1352 & ~n1355 ;
  assign n1363 = ~n1333 & n1362 ;
  assign n1365 = n1364 ^ n1363 ;
  assign n1366 = n1310 & n1365 ;
  assign n1371 = n1370 ^ n1366 ;
  assign n1218 = n672 & n999 ;
  assign n1221 = n1220 ^ n1218 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1226 = n1225 ^ n1223 ;
  assign n1209 = n972 & ~n999 ;
  assign n1212 = n1211 ^ n1209 ;
  assign n1214 = n1213 ^ n1212 ;
  assign n1217 = n1216 ^ n1214 ;
  assign n1227 = n1226 ^ n1217 ;
  assign n1207 = n584 & ~n666 ;
  assign n1206 = x40 & n666 ;
  assign n1208 = n1207 ^ n1206 ;
  assign n1228 = n1227 ^ n1208 ;
  assign n1241 = n995 & n999 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1246 = n1245 ^ n1244 ;
  assign n1249 = n1248 ^ n1246 ;
  assign n1232 = n992 & ~n999 ;
  assign n1235 = n1234 ^ n1232 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1240 = n1239 ^ n1237 ;
  assign n1250 = n1249 ^ n1240 ;
  assign n1230 = n588 & ~n666 ;
  assign n1229 = x41 & n666 ;
  assign n1231 = n1230 ^ n1229 ;
  assign n1251 = n1250 ^ n1231 ;
  assign n1252 = ~n1228 & ~n1251 ;
  assign n1169 = n999 & n1022 ;
  assign n1172 = n1171 ^ n1169 ;
  assign n1174 = n1173 ^ n1172 ;
  assign n1177 = n1176 ^ n1174 ;
  assign n1019 = ~n999 & n1018 ;
  assign n1054 = n1053 ^ n1019 ;
  assign n1155 = n1154 ^ n1054 ;
  assign n1168 = n1167 ^ n1155 ;
  assign n1178 = n1177 ^ n1168 ;
  assign n668 = n593 & ~n666 ;
  assign n667 = x42 & n666 ;
  assign n669 = n668 ^ n667 ;
  assign n1179 = n1178 ^ n669 ;
  assign n1192 = n999 & n1026 ;
  assign n1195 = n1194 ^ n1192 ;
  assign n1197 = n1196 ^ n1195 ;
  assign n1200 = n1199 ^ n1197 ;
  assign n1183 = ~n999 & n1045 ;
  assign n1186 = n1185 ^ n1183 ;
  assign n1188 = n1187 ^ n1186 ;
  assign n1191 = n1190 ^ n1188 ;
  assign n1201 = n1200 ^ n1191 ;
  assign n1181 = n597 & ~n666 ;
  assign n1180 = x43 & n666 ;
  assign n1182 = n1181 ^ n1180 ;
  assign n1261 = n1201 ^ n1182 ;
  assign n1262 = ~n1179 & ~n1261 ;
  assign n1263 = n1252 & n1262 ;
  assign n1891 = n1263 & n1282 ;
  assign n1892 = n1371 & n1891 ;
  assign n1356 = n1355 ^ n1352 ;
  assign n1357 = ~n1333 & ~n1356 ;
  assign n1358 = n1310 & n1357 ;
  assign n1359 = n1263 & n1358 ;
  assign n1889 = n1282 & ~n1359 ;
  assign n1257 = ~n1208 & n1227 ;
  assign n1255 = ~n1231 & n1250 ;
  assign n1256 = ~n1228 & n1255 ;
  assign n1258 = n1257 ^ n1256 ;
  assign n1887 = n1258 & n1282 ;
  assign n1204 = ~n669 & n1178 ;
  assign n1202 = ~n1182 & n1201 ;
  assign n1203 = ~n1179 & n1202 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1885 = n1252 & n1282 ;
  assign n1886 = n1205 & n1885 ;
  assign n1888 = n1887 ^ n1886 ;
  assign n1890 = n1889 ^ n1888 ;
  assign n1893 = n1892 ^ n1890 ;
  assign n1882 = n1263 & n1285 ;
  assign n1883 = n1371 & n1882 ;
  assign n1880 = n1285 & ~n1359 ;
  assign n1878 = ~n1258 & n1285 ;
  assign n1876 = n1252 & n1285 ;
  assign n1877 = n1205 & n1876 ;
  assign n1879 = n1878 ^ n1877 ;
  assign n1881 = n1880 ^ n1879 ;
  assign n1884 = n1883 ^ n1881 ;
  assign n1894 = n1893 ^ n1884 ;
  assign n2026 = n1875 & ~n1894 ;
  assign n1895 = n1894 ^ n1875 ;
  assign n1907 = n1638 & n1665 ;
  assign n1908 = n1907 ^ n1906 ;
  assign n1910 = n1909 ^ n1908 ;
  assign n1913 = n1912 ^ n1910 ;
  assign n1898 = ~n1638 & n1668 ;
  assign n1899 = n1898 ^ n1897 ;
  assign n1901 = n1900 ^ n1899 ;
  assign n1904 = n1903 ^ n1901 ;
  assign n1914 = n1913 ^ n1904 ;
  assign n1930 = n1263 & n1305 ;
  assign n1931 = n1371 & n1930 ;
  assign n1928 = n1305 & ~n1359 ;
  assign n1926 = n1258 & n1305 ;
  assign n1924 = n1252 & n1305 ;
  assign n1925 = n1205 & n1924 ;
  assign n1927 = n1926 ^ n1925 ;
  assign n1929 = n1928 ^ n1927 ;
  assign n1932 = n1931 ^ n1929 ;
  assign n1921 = n1263 & n1308 ;
  assign n1922 = n1371 & n1921 ;
  assign n1919 = n1308 & ~n1359 ;
  assign n1917 = ~n1258 & n1308 ;
  assign n1915 = n1252 & n1308 ;
  assign n1916 = n1205 & n1915 ;
  assign n1918 = n1917 ^ n1916 ;
  assign n1920 = n1919 ^ n1918 ;
  assign n1923 = n1922 ^ n1920 ;
  assign n1933 = n1932 ^ n1923 ;
  assign n2024 = n1914 & ~n1933 ;
  assign n2025 = ~n1895 & n2024 ;
  assign n2027 = n2026 ^ n2025 ;
  assign n1934 = n1933 ^ n1914 ;
  assign n1935 = ~n1895 & ~n1934 ;
  assign n1947 = n1638 & n1679 ;
  assign n1948 = n1947 ^ n1946 ;
  assign n1950 = n1949 ^ n1948 ;
  assign n1953 = n1952 ^ n1950 ;
  assign n1938 = ~n1638 & n1682 ;
  assign n1939 = n1938 ^ n1937 ;
  assign n1941 = n1940 ^ n1939 ;
  assign n1944 = n1943 ^ n1941 ;
  assign n1954 = n1953 ^ n1944 ;
  assign n1970 = n1263 & n1329 ;
  assign n1971 = n1371 & n1970 ;
  assign n1968 = n1329 & ~n1359 ;
  assign n1966 = n1258 & n1329 ;
  assign n1964 = n1252 & n1329 ;
  assign n1965 = n1205 & n1964 ;
  assign n1967 = n1966 ^ n1965 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n1972 = n1971 ^ n1969 ;
  assign n1961 = n1263 & n1332 ;
  assign n1962 = n1371 & n1961 ;
  assign n1959 = n1332 & ~n1359 ;
  assign n1957 = ~n1258 & n1332 ;
  assign n1955 = n1252 & n1332 ;
  assign n1956 = n1205 & n1955 ;
  assign n1958 = n1957 ^ n1956 ;
  assign n1960 = n1959 ^ n1958 ;
  assign n1963 = n1962 ^ n1960 ;
  assign n1973 = n1972 ^ n1963 ;
  assign n2021 = n1954 & ~n1973 ;
  assign n1974 = n1973 ^ n1954 ;
  assign n1986 = n1638 & n1695 ;
  assign n1987 = n1986 ^ n1985 ;
  assign n1989 = n1988 ^ n1987 ;
  assign n1992 = n1991 ^ n1989 ;
  assign n1977 = ~n1638 & n1686 ;
  assign n1978 = n1977 ^ n1976 ;
  assign n1980 = n1979 ^ n1978 ;
  assign n1983 = n1982 ^ n1980 ;
  assign n1993 = n1992 ^ n1983 ;
  assign n2009 = n1263 & n1352 ;
  assign n2010 = n1371 & n2009 ;
  assign n2007 = n1352 & ~n1359 ;
  assign n2005 = n1258 & n1352 ;
  assign n2003 = n1252 & n1352 ;
  assign n2004 = n1205 & n2003 ;
  assign n2006 = n2005 ^ n2004 ;
  assign n2008 = n2007 ^ n2006 ;
  assign n2011 = n2010 ^ n2008 ;
  assign n2000 = n1263 & n1355 ;
  assign n2001 = n1371 & n2000 ;
  assign n1998 = n1355 & ~n1359 ;
  assign n1996 = ~n1258 & n1355 ;
  assign n1994 = n1252 & n1355 ;
  assign n1995 = n1205 & n1994 ;
  assign n1997 = n1996 ^ n1995 ;
  assign n1999 = n1998 ^ n1997 ;
  assign n2002 = n2001 ^ n1999 ;
  assign n2012 = n2011 ^ n2002 ;
  assign n2019 = n1993 & ~n2012 ;
  assign n2020 = ~n1974 & n2019 ;
  assign n2022 = n2021 ^ n2020 ;
  assign n2023 = n1935 & n2022 ;
  assign n2028 = n2027 ^ n2023 ;
  assign n1717 = n1617 & n1638 ;
  assign n1718 = n1717 ^ n1716 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1723 = n1722 ^ n1720 ;
  assign n1639 = n1608 & ~n1638 ;
  assign n1640 = n1639 ^ n1634 ;
  assign n1701 = n1700 ^ n1640 ;
  assign n1714 = n1713 ^ n1701 ;
  assign n1724 = n1723 ^ n1714 ;
  assign n1381 = n1227 & n1263 ;
  assign n1382 = n1371 & n1381 ;
  assign n1379 = n1227 & ~n1359 ;
  assign n1377 = n1227 & n1258 ;
  assign n1375 = n1227 & n1252 ;
  assign n1376 = n1205 & n1375 ;
  assign n1378 = n1377 ^ n1376 ;
  assign n1380 = n1379 ^ n1378 ;
  assign n1383 = n1382 ^ n1380 ;
  assign n1372 = n1208 & n1263 ;
  assign n1373 = n1371 & n1372 ;
  assign n1360 = n1208 & ~n1359 ;
  assign n1259 = n1208 & ~n1258 ;
  assign n1253 = n1208 & n1252 ;
  assign n1254 = n1205 & n1253 ;
  assign n1260 = n1259 ^ n1254 ;
  assign n1361 = n1360 ^ n1260 ;
  assign n1374 = n1373 ^ n1361 ;
  assign n1384 = n1383 ^ n1374 ;
  assign n1725 = n1724 ^ n1384 ;
  assign n1760 = n1250 & n1263 ;
  assign n1761 = n1371 & n1760 ;
  assign n1758 = n1250 & ~n1359 ;
  assign n1756 = n1250 & n1258 ;
  assign n1754 = n1250 & n1252 ;
  assign n1755 = n1205 & n1754 ;
  assign n1757 = n1756 ^ n1755 ;
  assign n1759 = n1758 ^ n1757 ;
  assign n1762 = n1761 ^ n1759 ;
  assign n1751 = n1231 & n1263 ;
  assign n1752 = n1371 & n1751 ;
  assign n1749 = n1231 & ~n1359 ;
  assign n1747 = n1231 & ~n1258 ;
  assign n1745 = n1231 & n1252 ;
  assign n1746 = n1205 & n1745 ;
  assign n1748 = n1747 ^ n1746 ;
  assign n1750 = n1749 ^ n1748 ;
  assign n1753 = n1752 ^ n1750 ;
  assign n1763 = n1762 ^ n1753 ;
  assign n1737 = n1627 & n1638 ;
  assign n1738 = n1737 ^ n1736 ;
  assign n1740 = n1739 ^ n1738 ;
  assign n1743 = n1742 ^ n1740 ;
  assign n1728 = n1630 & ~n1638 ;
  assign n1729 = n1728 ^ n1727 ;
  assign n1731 = n1730 ^ n1729 ;
  assign n1734 = n1733 ^ n1731 ;
  assign n1744 = n1743 ^ n1734 ;
  assign n1764 = n1763 ^ n1744 ;
  assign n1765 = ~n1725 & ~n1764 ;
  assign n1800 = n1178 & n1263 ;
  assign n1801 = n1371 & n1800 ;
  assign n1798 = n1178 & ~n1359 ;
  assign n1796 = n1178 & n1258 ;
  assign n1794 = n1178 & n1252 ;
  assign n1795 = n1205 & n1794 ;
  assign n1797 = n1796 ^ n1795 ;
  assign n1799 = n1798 ^ n1797 ;
  assign n1802 = n1801 ^ n1799 ;
  assign n1791 = n669 & n1263 ;
  assign n1792 = n1371 & n1791 ;
  assign n1789 = n669 & ~n1359 ;
  assign n1787 = n669 & ~n1258 ;
  assign n1785 = n669 & n1252 ;
  assign n1786 = n1205 & n1785 ;
  assign n1788 = n1787 ^ n1786 ;
  assign n1790 = n1789 ^ n1788 ;
  assign n1793 = n1792 ^ n1790 ;
  assign n1803 = n1802 ^ n1793 ;
  assign n1777 = n1588 & n1638 ;
  assign n1778 = n1777 ^ n1776 ;
  assign n1780 = n1779 ^ n1778 ;
  assign n1783 = n1782 ^ n1780 ;
  assign n1768 = n1579 & ~n1638 ;
  assign n1769 = n1768 ^ n1767 ;
  assign n1771 = n1770 ^ n1769 ;
  assign n1774 = n1773 ^ n1771 ;
  assign n1784 = n1783 ^ n1774 ;
  assign n1804 = n1803 ^ n1784 ;
  assign n1835 = n1601 & n1638 ;
  assign n1836 = n1835 ^ n1834 ;
  assign n1838 = n1837 ^ n1836 ;
  assign n1841 = n1840 ^ n1838 ;
  assign n1826 = n1592 & ~n1638 ;
  assign n1827 = n1826 ^ n1825 ;
  assign n1829 = n1828 ^ n1827 ;
  assign n1832 = n1831 ^ n1829 ;
  assign n1842 = n1841 ^ n1832 ;
  assign n1820 = n1201 & n1263 ;
  assign n1821 = n1371 & n1820 ;
  assign n1818 = n1201 & ~n1359 ;
  assign n1816 = n1201 & n1258 ;
  assign n1814 = n1201 & n1252 ;
  assign n1815 = n1205 & n1814 ;
  assign n1817 = n1816 ^ n1815 ;
  assign n1819 = n1818 ^ n1817 ;
  assign n1822 = n1821 ^ n1819 ;
  assign n1811 = n1182 & n1263 ;
  assign n1812 = n1371 & n1811 ;
  assign n1809 = n1182 & ~n1359 ;
  assign n1807 = n1182 & ~n1258 ;
  assign n1805 = n1182 & n1252 ;
  assign n1806 = n1205 & n1805 ;
  assign n1808 = n1807 ^ n1806 ;
  assign n1810 = n1809 ^ n1808 ;
  assign n1813 = n1812 ^ n1810 ;
  assign n1823 = n1822 ^ n1813 ;
  assign n1854 = n1842 ^ n1823 ;
  assign n1855 = ~n1804 & ~n1854 ;
  assign n1856 = n1765 & n1855 ;
  assign n2312 = n1856 & n1875 ;
  assign n2313 = n2028 & n2312 ;
  assign n2013 = n2012 ^ n1993 ;
  assign n2014 = ~n1974 & ~n2013 ;
  assign n2015 = n1935 & n2014 ;
  assign n2016 = n1856 & n2015 ;
  assign n2310 = n1875 & ~n2016 ;
  assign n1850 = ~n1384 & n1724 ;
  assign n1848 = n1744 & ~n1763 ;
  assign n1849 = ~n1725 & n1848 ;
  assign n1851 = n1850 ^ n1849 ;
  assign n1845 = n1784 & ~n1803 ;
  assign n1843 = ~n1823 & n1842 ;
  assign n1844 = ~n1804 & n1843 ;
  assign n1846 = n1845 ^ n1844 ;
  assign n1847 = n1765 & n1846 ;
  assign n1852 = n1851 ^ n1847 ;
  assign n2309 = n1852 & n1875 ;
  assign n2311 = n2310 ^ n2309 ;
  assign n2314 = n2313 ^ n2311 ;
  assign n2306 = n1856 & n1894 ;
  assign n2307 = n2028 & n2306 ;
  assign n2304 = n1894 & ~n2016 ;
  assign n2303 = ~n1852 & n1894 ;
  assign n2305 = n2304 ^ n2303 ;
  assign n2308 = n2307 ^ n2305 ;
  assign n2315 = n2314 ^ n2308 ;
  assign n2387 = n2302 & ~n2315 ;
  assign n2316 = n2315 ^ n2302 ;
  assign n2318 = n2118 & ~n2230 ;
  assign n2317 = n2109 & n2230 ;
  assign n2319 = n2318 ^ n2317 ;
  assign n2329 = n1856 & n1914 ;
  assign n2330 = n2028 & n2329 ;
  assign n2327 = n1914 & ~n2016 ;
  assign n2326 = n1852 & n1914 ;
  assign n2328 = n2327 ^ n2326 ;
  assign n2331 = n2330 ^ n2328 ;
  assign n2323 = n1856 & n1933 ;
  assign n2324 = n2028 & n2323 ;
  assign n2321 = n1933 & ~n2016 ;
  assign n2320 = ~n1852 & n1933 ;
  assign n2322 = n2321 ^ n2320 ;
  assign n2325 = n2324 ^ n2322 ;
  assign n2332 = n2331 ^ n2325 ;
  assign n2385 = n2319 & ~n2332 ;
  assign n2386 = ~n2316 & n2385 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2333 = n2332 ^ n2319 ;
  assign n2334 = ~n2316 & ~n2333 ;
  assign n2336 = n2129 & ~n2230 ;
  assign n2335 = n2132 & n2230 ;
  assign n2337 = n2336 ^ n2335 ;
  assign n2347 = n1856 & n1954 ;
  assign n2348 = n2028 & n2347 ;
  assign n2345 = n1954 & ~n2016 ;
  assign n2344 = n1852 & n1954 ;
  assign n2346 = n2345 ^ n2344 ;
  assign n2349 = n2348 ^ n2346 ;
  assign n2341 = n1856 & n1973 ;
  assign n2342 = n2028 & n2341 ;
  assign n2339 = n1973 & ~n2016 ;
  assign n2338 = ~n1852 & n1973 ;
  assign n2340 = n2339 ^ n2338 ;
  assign n2343 = n2342 ^ n2340 ;
  assign n2350 = n2349 ^ n2343 ;
  assign n2382 = n2337 & ~n2350 ;
  assign n2351 = n2350 ^ n2337 ;
  assign n2353 = n2142 & ~n2230 ;
  assign n2352 = n2145 & n2230 ;
  assign n2354 = n2353 ^ n2352 ;
  assign n2370 = n1856 & n1993 ;
  assign n2371 = n2028 & n2370 ;
  assign n2368 = n1993 & ~n2016 ;
  assign n2366 = n1851 & n1993 ;
  assign n2364 = n1765 & n1993 ;
  assign n2365 = n1846 & n2364 ;
  assign n2367 = n2366 ^ n2365 ;
  assign n2369 = n2368 ^ n2367 ;
  assign n2372 = n2371 ^ n2369 ;
  assign n2361 = n1856 & n2012 ;
  assign n2362 = n2028 & n2361 ;
  assign n2359 = n2012 & ~n2016 ;
  assign n2357 = ~n1851 & n2012 ;
  assign n2355 = n1765 & n2012 ;
  assign n2356 = n1846 & n2355 ;
  assign n2358 = n2357 ^ n2356 ;
  assign n2360 = n2359 ^ n2358 ;
  assign n2363 = n2362 ^ n2360 ;
  assign n2373 = n2372 ^ n2363 ;
  assign n2380 = n2354 & ~n2373 ;
  assign n2381 = ~n2351 & n2380 ;
  assign n2383 = n2382 ^ n2381 ;
  assign n2384 = n2334 & n2383 ;
  assign n2389 = n2388 ^ n2384 ;
  assign n2232 = n2050 & ~n2230 ;
  assign n2231 = n2041 & n2230 ;
  assign n2233 = n2232 ^ n2231 ;
  assign n2035 = n1724 & n1856 ;
  assign n2036 = n2028 & n2035 ;
  assign n2033 = n1724 & ~n2016 ;
  assign n2032 = n1724 & n1852 ;
  assign n2034 = n2033 ^ n2032 ;
  assign n2037 = n2036 ^ n2034 ;
  assign n2029 = n1384 & n1856 ;
  assign n2030 = n2028 & n2029 ;
  assign n2017 = n1384 & ~n2016 ;
  assign n1853 = n1384 & ~n1852 ;
  assign n2018 = n2017 ^ n1853 ;
  assign n2031 = n2030 ^ n2018 ;
  assign n2038 = n2037 ^ n2031 ;
  assign n2234 = n2233 ^ n2038 ;
  assign n2247 = n1744 & n1856 ;
  assign n2248 = n2028 & n2247 ;
  assign n2245 = n1744 & ~n2016 ;
  assign n2244 = n1744 & n1852 ;
  assign n2246 = n2245 ^ n2244 ;
  assign n2249 = n2248 ^ n2246 ;
  assign n2241 = n1763 & n1856 ;
  assign n2242 = n2028 & n2241 ;
  assign n2239 = n1763 & ~n2016 ;
  assign n2238 = n1763 & ~n1852 ;
  assign n2240 = n2239 ^ n2238 ;
  assign n2243 = n2242 ^ n2240 ;
  assign n2250 = n2249 ^ n2243 ;
  assign n2236 = n2060 & ~n2230 ;
  assign n2235 = n2063 & n2230 ;
  assign n2237 = n2236 ^ n2235 ;
  assign n2251 = n2250 ^ n2237 ;
  assign n2252 = ~n2234 & ~n2251 ;
  assign n2265 = n1784 & n1856 ;
  assign n2266 = n2028 & n2265 ;
  assign n2263 = n1784 & ~n2016 ;
  assign n2262 = n1784 & n1852 ;
  assign n2264 = n2263 ^ n2262 ;
  assign n2267 = n2266 ^ n2264 ;
  assign n2259 = n1803 & n1856 ;
  assign n2260 = n2028 & n2259 ;
  assign n2257 = n1803 & ~n2016 ;
  assign n2256 = n1803 & ~n1852 ;
  assign n2258 = n2257 ^ n2256 ;
  assign n2261 = n2260 ^ n2258 ;
  assign n2268 = n2267 ^ n2261 ;
  assign n2254 = n2077 & ~n2230 ;
  assign n2253 = n2068 & n2230 ;
  assign n2255 = n2254 ^ n2253 ;
  assign n2269 = n2268 ^ n2255 ;
  assign n2284 = n2090 & ~n2230 ;
  assign n2283 = n2081 & n2230 ;
  assign n2285 = n2284 ^ n2283 ;
  assign n2279 = n1842 & n1856 ;
  assign n2280 = n2028 & n2279 ;
  assign n2277 = n1842 & ~n2016 ;
  assign n2276 = n1842 & n1852 ;
  assign n2278 = n2277 ^ n2276 ;
  assign n2281 = n2280 ^ n2278 ;
  assign n2273 = n1823 & n1856 ;
  assign n2274 = n2028 & n2273 ;
  assign n2271 = n1823 & ~n2016 ;
  assign n2270 = n1823 & ~n1852 ;
  assign n2272 = n2271 ^ n2270 ;
  assign n2275 = n2274 ^ n2272 ;
  assign n2282 = n2281 ^ n2275 ;
  assign n2297 = n2285 ^ n2282 ;
  assign n2298 = ~n2269 & ~n2297 ;
  assign n2299 = n2252 & n2298 ;
  assign n2396 = n2233 & n2299 ;
  assign n2397 = n2389 & n2396 ;
  assign n2374 = n2373 ^ n2354 ;
  assign n2375 = ~n2351 & ~n2374 ;
  assign n2376 = n2334 & n2375 ;
  assign n2377 = n2299 & n2376 ;
  assign n2394 = n2233 & ~n2377 ;
  assign n2293 = ~n2038 & n2233 ;
  assign n2291 = n2237 & ~n2250 ;
  assign n2292 = ~n2234 & n2291 ;
  assign n2294 = n2293 ^ n2292 ;
  assign n2288 = n2255 & ~n2268 ;
  assign n2286 = ~n2282 & n2285 ;
  assign n2287 = ~n2269 & n2286 ;
  assign n2289 = n2288 ^ n2287 ;
  assign n2290 = n2252 & n2289 ;
  assign n2295 = n2294 ^ n2290 ;
  assign n2393 = n2233 & n2295 ;
  assign n2395 = n2394 ^ n2393 ;
  assign n2398 = n2397 ^ n2395 ;
  assign n2390 = n2038 & n2299 ;
  assign n2391 = n2389 & n2390 ;
  assign n2378 = n2038 & ~n2377 ;
  assign n2296 = n2038 & ~n2295 ;
  assign n2379 = n2378 ^ n2296 ;
  assign n2392 = n2391 ^ n2379 ;
  assign n2399 = n2398 ^ n2392 ;
  assign n2403 = n2402 ^ n2399 ;
  assign n2418 = n2063 & ~n2230 ;
  assign n2417 = n2060 & n2230 ;
  assign n2419 = n2418 ^ n2417 ;
  assign n2413 = n2237 & n2299 ;
  assign n2414 = n2389 & n2413 ;
  assign n2411 = n2237 & ~n2377 ;
  assign n2410 = n2237 & n2295 ;
  assign n2412 = n2411 ^ n2410 ;
  assign n2415 = n2414 ^ n2412 ;
  assign n2407 = n2250 & n2299 ;
  assign n2408 = n2389 & n2407 ;
  assign n2405 = n2250 & ~n2377 ;
  assign n2404 = n2250 & ~n2295 ;
  assign n2406 = n2405 ^ n2404 ;
  assign n2409 = n2408 ^ n2406 ;
  assign n2416 = n2415 ^ n2409 ;
  assign n2420 = n2419 ^ n2416 ;
  assign n2421 = ~n2403 & ~n2420 ;
  assign n2423 = n2068 & ~n2230 ;
  assign n2422 = n2077 & n2230 ;
  assign n2424 = n2423 ^ n2422 ;
  assign n2434 = n2255 & n2299 ;
  assign n2435 = n2389 & n2434 ;
  assign n2432 = n2255 & ~n2377 ;
  assign n2431 = n2255 & n2295 ;
  assign n2433 = n2432 ^ n2431 ;
  assign n2436 = n2435 ^ n2433 ;
  assign n2428 = n2268 & n2299 ;
  assign n2429 = n2389 & n2428 ;
  assign n2426 = n2268 & ~n2377 ;
  assign n2425 = n2268 & ~n2295 ;
  assign n2427 = n2426 ^ n2425 ;
  assign n2430 = n2429 ^ n2427 ;
  assign n2437 = n2436 ^ n2430 ;
  assign n2573 = n2424 & ~n2437 ;
  assign n2438 = n2437 ^ n2424 ;
  assign n2530 = n2299 & n2389 ;
  assign n2531 = n2530 ^ n2295 ;
  assign n2532 = n2531 ^ n2377 ;
  assign n2453 = n2081 & ~n2230 ;
  assign n2452 = n2090 & n2230 ;
  assign n2454 = n2453 ^ n2452 ;
  assign n2569 = ~n2282 & n2454 ;
  assign n2570 = n2532 & n2569 ;
  assign n2567 = ~n2285 & n2454 ;
  assign n2568 = ~n2532 & n2567 ;
  assign n2571 = n2570 ^ n2568 ;
  assign n2572 = ~n2438 & n2571 ;
  assign n2574 = n2573 ^ n2572 ;
  assign n2575 = n2421 & n2574 ;
  assign n2565 = ~n2399 & n2402 ;
  assign n2563 = ~n2403 & n2419 ;
  assign n2564 = ~n2416 & n2563 ;
  assign n2566 = n2565 ^ n2564 ;
  assign n2576 = n2575 ^ n2566 ;
  assign n2448 = n2285 & n2299 ;
  assign n2449 = n2389 & n2448 ;
  assign n2446 = n2285 & ~n2377 ;
  assign n2445 = n2285 & n2295 ;
  assign n2447 = n2446 ^ n2445 ;
  assign n2450 = n2449 ^ n2447 ;
  assign n2442 = n2282 & n2299 ;
  assign n2443 = n2389 & n2442 ;
  assign n2440 = n2282 & ~n2377 ;
  assign n2439 = n2282 & ~n2295 ;
  assign n2441 = n2440 ^ n2439 ;
  assign n2444 = n2443 ^ n2441 ;
  assign n2451 = n2450 ^ n2444 ;
  assign n2455 = n2454 ^ n2451 ;
  assign n2456 = ~n2438 & ~n2455 ;
  assign n2457 = n2421 & n2456 ;
  assign n2459 = n2096 & ~n2230 ;
  assign n2458 = n2105 & n2230 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2470 = n2299 & n2302 ;
  assign n2471 = n2389 & n2470 ;
  assign n2468 = n2302 & ~n2377 ;
  assign n2467 = n2295 & n2302 ;
  assign n2469 = n2468 ^ n2467 ;
  assign n2472 = n2471 ^ n2469 ;
  assign n2464 = n2299 & n2315 ;
  assign n2465 = n2389 & n2464 ;
  assign n2462 = n2315 & ~n2377 ;
  assign n2461 = ~n2295 & n2315 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2466 = n2465 ^ n2463 ;
  assign n2473 = n2472 ^ n2466 ;
  assign n2559 = n2460 & ~n2473 ;
  assign n2474 = n2473 ^ n2460 ;
  assign n2489 = n2109 & ~n2230 ;
  assign n2488 = n2118 & n2230 ;
  assign n2490 = n2489 ^ n2488 ;
  assign n2555 = ~n2332 & n2490 ;
  assign n2556 = n2532 & n2555 ;
  assign n2553 = ~n2319 & n2490 ;
  assign n2554 = ~n2532 & n2553 ;
  assign n2557 = n2556 ^ n2554 ;
  assign n2558 = ~n2474 & n2557 ;
  assign n2560 = n2559 ^ n2558 ;
  assign n2484 = n2299 & n2319 ;
  assign n2485 = n2389 & n2484 ;
  assign n2482 = n2319 & ~n2377 ;
  assign n2481 = n2295 & n2319 ;
  assign n2483 = n2482 ^ n2481 ;
  assign n2486 = n2485 ^ n2483 ;
  assign n2478 = n2299 & n2332 ;
  assign n2479 = n2389 & n2478 ;
  assign n2476 = n2332 & ~n2377 ;
  assign n2475 = ~n2295 & n2332 ;
  assign n2477 = n2476 ^ n2475 ;
  assign n2480 = n2479 ^ n2477 ;
  assign n2487 = n2486 ^ n2480 ;
  assign n2491 = n2490 ^ n2487 ;
  assign n2492 = ~n2474 & ~n2491 ;
  assign n2507 = n2132 & ~n2230 ;
  assign n2506 = n2129 & n2230 ;
  assign n2508 = n2507 ^ n2506 ;
  assign n2549 = ~n2337 & n2508 ;
  assign n2550 = ~n2532 & n2549 ;
  assign n2524 = n2145 & ~n2230 ;
  assign n2523 = n2142 & n2230 ;
  assign n2525 = n2524 ^ n2523 ;
  assign n2538 = ~n2354 & n2525 ;
  assign n2544 = n2508 & n2538 ;
  assign n2545 = ~n2532 & n2544 ;
  assign n2535 = ~n2373 & n2525 ;
  assign n2542 = n2508 & n2535 ;
  assign n2543 = n2532 & n2542 ;
  assign n2546 = n2545 ^ n2543 ;
  assign n2539 = ~n2337 & n2538 ;
  assign n2540 = ~n2532 & n2539 ;
  assign n2536 = ~n2350 & n2535 ;
  assign n2537 = n2532 & n2536 ;
  assign n2541 = n2540 ^ n2537 ;
  assign n2547 = n2546 ^ n2541 ;
  assign n2533 = ~n2350 & n2508 ;
  assign n2534 = n2532 & n2533 ;
  assign n2548 = n2547 ^ n2534 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2552 = n2492 & n2551 ;
  assign n2561 = n2560 ^ n2552 ;
  assign n2562 = n2457 & n2561 ;
  assign n2577 = n2576 ^ n2562 ;
  assign n2502 = n2299 & n2337 ;
  assign n2503 = n2389 & n2502 ;
  assign n2500 = n2337 & ~n2377 ;
  assign n2499 = n2295 & n2337 ;
  assign n2501 = n2500 ^ n2499 ;
  assign n2504 = n2503 ^ n2501 ;
  assign n2496 = n2299 & n2350 ;
  assign n2497 = n2389 & n2496 ;
  assign n2494 = n2350 & ~n2377 ;
  assign n2493 = ~n2295 & n2350 ;
  assign n2495 = n2494 ^ n2493 ;
  assign n2498 = n2497 ^ n2495 ;
  assign n2505 = n2504 ^ n2498 ;
  assign n2509 = n2508 ^ n2505 ;
  assign n2519 = n2299 & n2354 ;
  assign n2520 = n2389 & n2519 ;
  assign n2517 = n2354 & ~n2377 ;
  assign n2516 = n2295 & n2354 ;
  assign n2518 = n2517 ^ n2516 ;
  assign n2521 = n2520 ^ n2518 ;
  assign n2513 = n2299 & n2373 ;
  assign n2514 = n2389 & n2513 ;
  assign n2511 = n2373 & ~n2377 ;
  assign n2510 = ~n2295 & n2373 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2515 = n2514 ^ n2512 ;
  assign n2522 = n2521 ^ n2515 ;
  assign n2526 = n2525 ^ n2522 ;
  assign n2527 = ~n2509 & ~n2526 ;
  assign n2528 = n2492 & n2527 ;
  assign n2529 = n2457 & n2528 ;
  assign n2578 = n2577 ^ n2529 ;
  assign n2580 = n2402 & ~n2578 ;
  assign n2579 = n2399 & n2578 ;
  assign n2581 = n2580 ^ n2579 ;
  assign n2583 = n2419 & ~n2578 ;
  assign n2582 = n2416 & n2578 ;
  assign n2584 = n2583 ^ n2582 ;
  assign n2586 = n2424 & ~n2578 ;
  assign n2585 = n2437 & n2578 ;
  assign n2587 = n2586 ^ n2585 ;
  assign n2589 = n2454 & ~n2578 ;
  assign n2588 = n2451 & n2578 ;
  assign n2590 = n2589 ^ n2588 ;
  assign n2592 = n2460 & ~n2578 ;
  assign n2591 = n2473 & n2578 ;
  assign n2593 = n2592 ^ n2591 ;
  assign n2595 = n2490 & ~n2578 ;
  assign n2594 = n2487 & n2578 ;
  assign n2596 = n2595 ^ n2594 ;
  assign n2598 = n2508 & ~n2578 ;
  assign n2597 = n2505 & n2578 ;
  assign n2599 = n2598 ^ n2597 ;
  assign n2601 = n2525 & ~n2578 ;
  assign n2600 = n2522 & n2578 ;
  assign n2602 = n2601 ^ n2600 ;
  assign n2604 = n2399 & ~n2578 ;
  assign n2603 = n2402 & n2578 ;
  assign n2605 = n2604 ^ n2603 ;
  assign n2607 = n2416 & ~n2578 ;
  assign n2606 = n2419 & n2578 ;
  assign n2608 = n2607 ^ n2606 ;
  assign n2610 = n2437 & ~n2578 ;
  assign n2609 = n2424 & n2578 ;
  assign n2611 = n2610 ^ n2609 ;
  assign n2613 = n2451 & ~n2578 ;
  assign n2612 = n2454 & n2578 ;
  assign n2614 = n2613 ^ n2612 ;
  assign n2616 = n2473 & ~n2578 ;
  assign n2615 = n2460 & n2578 ;
  assign n2617 = n2616 ^ n2615 ;
  assign n2619 = n2487 & ~n2578 ;
  assign n2618 = n2490 & n2578 ;
  assign n2620 = n2619 ^ n2618 ;
  assign n2622 = n2505 & ~n2578 ;
  assign n2621 = n2508 & n2578 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2625 = n2522 & ~n2578 ;
  assign n2624 = n2525 & n2578 ;
  assign n2626 = n2625 ^ n2624 ;
  assign n2628 = n2038 & ~n2532 ;
  assign n2627 = n2233 & n2532 ;
  assign n2629 = n2628 ^ n2627 ;
  assign n2631 = n2250 & ~n2532 ;
  assign n2630 = n2237 & n2532 ;
  assign n2632 = n2631 ^ n2630 ;
  assign n2634 = n2268 & ~n2532 ;
  assign n2633 = n2255 & n2532 ;
  assign n2635 = n2634 ^ n2633 ;
  assign n2637 = n2282 & ~n2532 ;
  assign n2636 = n2285 & n2532 ;
  assign n2638 = n2637 ^ n2636 ;
  assign n2640 = n2315 & ~n2532 ;
  assign n2639 = n2302 & n2532 ;
  assign n2641 = n2640 ^ n2639 ;
  assign n2643 = n2332 & ~n2532 ;
  assign n2642 = n2319 & n2532 ;
  assign n2644 = n2643 ^ n2642 ;
  assign n2646 = n2350 & ~n2532 ;
  assign n2645 = n2337 & n2532 ;
  assign n2647 = n2646 ^ n2645 ;
  assign n2649 = n2373 & ~n2532 ;
  assign n2648 = n2354 & n2532 ;
  assign n2650 = n2649 ^ n2648 ;
  assign n2651 = n1856 & n2028 ;
  assign n2652 = n2651 ^ n1852 ;
  assign n2653 = n2652 ^ n2016 ;
  assign n2655 = n1384 & ~n2653 ;
  assign n2654 = n1724 & n2653 ;
  assign n2656 = n2655 ^ n2654 ;
  assign n2658 = n1763 & ~n2653 ;
  assign n2657 = n1744 & n2653 ;
  assign n2659 = n2658 ^ n2657 ;
  assign n2661 = n1803 & ~n2653 ;
  assign n2660 = n1784 & n2653 ;
  assign n2662 = n2661 ^ n2660 ;
  assign n2664 = n1823 & ~n2653 ;
  assign n2663 = n1842 & n2653 ;
  assign n2665 = n2664 ^ n2663 ;
  assign n2667 = n1894 & ~n2653 ;
  assign n2666 = n1875 & n2653 ;
  assign n2668 = n2667 ^ n2666 ;
  assign n2670 = n1933 & ~n2653 ;
  assign n2669 = n1914 & n2653 ;
  assign n2671 = n2670 ^ n2669 ;
  assign n2673 = n1973 & ~n2653 ;
  assign n2672 = n1954 & n2653 ;
  assign n2674 = n2673 ^ n2672 ;
  assign n2676 = n2012 & ~n2653 ;
  assign n2675 = n1993 & n2653 ;
  assign n2677 = n2676 ^ n2675 ;
  assign n2679 = n1205 & n1252 ;
  assign n2680 = n2679 ^ n1258 ;
  assign n2678 = n1263 & n1371 ;
  assign n2681 = n2680 ^ n2678 ;
  assign n2682 = n2681 ^ n1359 ;
  assign n2684 = n1208 & ~n2682 ;
  assign n2683 = n1227 & n2682 ;
  assign n2685 = n2684 ^ n2683 ;
  assign n2687 = n1231 & ~n2682 ;
  assign n2686 = n1250 & n2682 ;
  assign n2688 = n2687 ^ n2686 ;
  assign n2690 = n669 & ~n2682 ;
  assign n2689 = n1178 & n2682 ;
  assign n2691 = n2690 ^ n2689 ;
  assign n2693 = n1182 & ~n2682 ;
  assign n2692 = n1201 & n2682 ;
  assign n2694 = n2693 ^ n2692 ;
  assign n2696 = n1285 & ~n2682 ;
  assign n2695 = n1282 & n2682 ;
  assign n2697 = n2696 ^ n2695 ;
  assign n2699 = n1308 & ~n2682 ;
  assign n2698 = n1305 & n2682 ;
  assign n2700 = n2699 ^ n2698 ;
  assign n2702 = n1332 & ~n2682 ;
  assign n2701 = n1329 & n2682 ;
  assign n2703 = n2702 ^ n2701 ;
  assign n2705 = n1355 & ~n2682 ;
  assign n2704 = n1352 & n2682 ;
  assign n2706 = n2705 ^ n2704 ;
  assign n2708 = x40 & ~n666 ;
  assign n2707 = n584 & n666 ;
  assign n2709 = n2708 ^ n2707 ;
  assign n2711 = x41 & ~n666 ;
  assign n2710 = n588 & n666 ;
  assign n2712 = n2711 ^ n2710 ;
  assign n2714 = x42 & ~n666 ;
  assign n2713 = n593 & n666 ;
  assign n2715 = n2714 ^ n2713 ;
  assign n2717 = x43 & ~n666 ;
  assign n2716 = n597 & n666 ;
  assign n2718 = n2717 ^ n2716 ;
  assign n2720 = x44 & ~n666 ;
  assign n2719 = n603 & n666 ;
  assign n2721 = n2720 ^ n2719 ;
  assign n2723 = x45 & ~n666 ;
  assign n2722 = n607 & n666 ;
  assign n2724 = n2723 ^ n2722 ;
  assign n2726 = x46 & ~n666 ;
  assign n2725 = n612 & n666 ;
  assign n2727 = n2726 ^ n2725 ;
  assign n2729 = x47 & ~n666 ;
  assign n2728 = n616 & n666 ;
  assign n2730 = n2729 ^ n2728 ;
  assign y0 = n2581 ;
  assign y1 = n2584 ;
  assign y2 = n2587 ;
  assign y3 = n2590 ;
  assign y4 = n2593 ;
  assign y5 = n2596 ;
  assign y6 = n2599 ;
  assign y7 = n2602 ;
  assign y8 = n2605 ;
  assign y9 = n2608 ;
  assign y10 = n2611 ;
  assign y11 = n2614 ;
  assign y12 = n2617 ;
  assign y13 = n2620 ;
  assign y14 = n2623 ;
  assign y15 = n2626 ;
  assign y16 = n2629 ;
  assign y17 = n2632 ;
  assign y18 = n2635 ;
  assign y19 = n2638 ;
  assign y20 = n2641 ;
  assign y21 = n2644 ;
  assign y22 = n2647 ;
  assign y23 = n2650 ;
  assign y24 = n2656 ;
  assign y25 = n2659 ;
  assign y26 = n2662 ;
  assign y27 = n2665 ;
  assign y28 = n2668 ;
  assign y29 = n2671 ;
  assign y30 = n2674 ;
  assign y31 = n2677 ;
  assign y32 = n2685 ;
  assign y33 = n2688 ;
  assign y34 = n2691 ;
  assign y35 = n2694 ;
  assign y36 = n2697 ;
  assign y37 = n2700 ;
  assign y38 = n2703 ;
  assign y39 = n2706 ;
  assign y40 = n2709 ;
  assign y41 = n2712 ;
  assign y42 = n2715 ;
  assign y43 = n2718 ;
  assign y44 = n2721 ;
  assign y45 = n2724 ;
  assign y46 = n2727 ;
  assign y47 = n2730 ;
endmodule
