module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 ;
  assign n61 = x20 & x21 ;
  assign n62 = n61 ^ x20 ;
  assign n63 = x22 & x23 ;
  assign n64 = n63 ^ x23 ;
  assign n65 = ~x1 & ~x2 ;
  assign n66 = n64 & n65 ;
  assign n67 = n62 & n66 ;
  assign n68 = x9 & x10 ;
  assign n69 = n68 ^ x9 ;
  assign n70 = x7 & x8 ;
  assign n71 = n70 ^ x7 ;
  assign n72 = n71 ^ x8 ;
  assign n73 = n69 & ~n72 ;
  assign n74 = x3 & x4 ;
  assign n75 = n74 ^ x3 ;
  assign n76 = n75 ^ x4 ;
  assign n77 = x5 & x6 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = n78 ^ x6 ;
  assign n80 = ~n76 & ~n79 ;
  assign n81 = n73 & n80 ;
  assign n82 = x24 & x25 ;
  assign n83 = x26 & n82 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = x13 & x14 ;
  assign n86 = n85 ^ x14 ;
  assign n87 = x18 & x19 ;
  assign n88 = n87 ^ x19 ;
  assign n89 = n86 & n88 ;
  assign n90 = n84 & n89 ;
  assign n91 = n81 & n90 ;
  assign n92 = n67 & n91 ;
  assign n93 = n69 ^ x10 ;
  assign n94 = x11 & n93 ;
  assign n95 = x12 & x13 ;
  assign n96 = n95 ^ x12 ;
  assign n97 = n96 ^ x13 ;
  assign n98 = x14 & x15 ;
  assign n99 = n97 & n98 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = n94 & n100 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = n102 ^ n98 ;
  assign n104 = x16 & n103 ;
  assign n105 = ~x12 & n94 ;
  assign n106 = ~x11 & x12 ;
  assign n107 = ~n93 & n106 ;
  assign n108 = ~n105 & ~n107 ;
  assign n109 = ~n104 & ~n108 ;
  assign n110 = n92 & n109 ;
  assign n122 = x23 & x24 ;
  assign n128 = x25 & n122 ;
  assign n115 = ~x16 & x17 ;
  assign n111 = x19 & x20 ;
  assign n116 = x18 & n111 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n115 & n117 ;
  assign n119 = n103 & n118 ;
  assign n120 = n119 ^ n118 ;
  assign n112 = ~x17 & ~x18 ;
  assign n113 = n111 & n112 ;
  assign n114 = n113 ^ n111 ;
  assign n121 = n120 ^ n114 ;
  assign n123 = ~x21 & ~x22 ;
  assign n124 = x25 & n123 ;
  assign n125 = n122 & n124 ;
  assign n126 = n121 & n125 ;
  assign n127 = n126 ^ n125 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = x27 & x28 ;
  assign n131 = x29 & n130 ;
  assign n132 = ~x26 & n131 ;
  assign n133 = n129 & n132 ;
  assign n134 = n133 ^ n132 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = ~n103 & n115 ;
  assign n137 = n136 ^ x17 ;
  assign n138 = x14 & ~n97 ;
  assign n139 = ~n94 & n138 ;
  assign n140 = n139 ^ x14 ;
  assign n141 = n140 ^ x15 ;
  assign n142 = n137 & ~n141 ;
  assign n143 = n135 & n142 ;
  assign n144 = n110 & n143 ;
  assign n145 = n144 ^ n135 ;
  assign n146 = x19 & x25 ;
  assign n147 = x26 & n146 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = x15 & x16 ;
  assign n150 = n149 ^ x15 ;
  assign n151 = n97 & n150 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n148 & n152 ;
  assign n154 = n131 & n153 ;
  assign n155 = n62 & n64 ;
  assign n156 = x0 & x1 ;
  assign n157 = n93 & n156 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n155 & n158 ;
  assign n160 = x6 & x7 ;
  assign n161 = x8 & x11 ;
  assign n162 = n160 & n161 ;
  assign n163 = x2 & x3 ;
  assign n164 = x4 & x5 ;
  assign n165 = n163 & n164 ;
  assign n166 = n162 & n165 ;
  assign n167 = n159 & n166 ;
  assign n168 = n154 & n167 ;
  assign n172 = ~n94 & ~n97 ;
  assign n173 = n172 ^ x14 ;
  assign n180 = n168 & n173 ;
  assign n181 = n180 ^ n168 ;
  assign n169 = ~x16 & ~x17 ;
  assign n170 = ~n103 & n169 ;
  assign n171 = n170 ^ n168 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = n173 & ~n174 ;
  assign n176 = n175 ^ n170 ;
  assign n177 = n171 & ~n176 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n178 ^ n168 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = ~x18 & n115 ;
  assign n184 = ~n103 & n183 ;
  assign n185 = n184 ^ n112 ;
  assign n195 = ~x24 & n185 ;
  assign n196 = n135 & n195 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n182 & n197 ;
  assign n186 = x23 & n123 ;
  assign n187 = n121 & n186 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = n188 ^ x23 ;
  assign n190 = n185 & n189 ;
  assign n191 = n190 ^ n185 ;
  assign n192 = n135 & n191 ;
  assign n193 = n192 ^ n191 ;
  assign n194 = n182 & n193 ;
  assign n199 = n198 ^ n194 ;
  assign n200 = n199 ^ n135 ;
  assign n201 = n145 & n200 ;
  assign n202 = n201 ^ n200 ;
  assign n399 = n181 ^ n170 ;
  assign n400 = n185 ^ n170 ;
  assign n401 = n185 & n400 ;
  assign n402 = n401 ^ n185 ;
  assign n403 = n402 ^ n400 ;
  assign n404 = n403 ^ n170 ;
  assign n405 = n399 & ~n404 ;
  assign n406 = n405 ^ n404 ;
  assign n407 = n406 ^ n403 ;
  assign n408 = n407 ^ n181 ;
  assign n409 = x23 & ~n121 ;
  assign n410 = n123 & n409 ;
  assign n411 = n410 ^ x23 ;
  assign n412 = n411 ^ x24 ;
  assign n413 = n408 & n412 ;
  assign n217 = x45 & x46 ;
  assign n218 = n217 ^ x45 ;
  assign n224 = x44 & n218 ;
  assign n210 = x39 & x40 ;
  assign n211 = n210 ^ x39 ;
  assign n212 = n211 ^ x40 ;
  assign n213 = x41 & x42 ;
  assign n214 = n213 ^ x41 ;
  assign n215 = n212 & n214 ;
  assign n216 = n215 ^ x42 ;
  assign n219 = x43 & x44 ;
  assign n220 = n219 ^ x44 ;
  assign n221 = n218 & n220 ;
  assign n222 = n216 & n221 ;
  assign n223 = n222 ^ n221 ;
  assign n225 = n224 ^ n223 ;
  assign n226 = n225 ^ x46 ;
  assign n203 = x49 & x50 ;
  assign n204 = x52 & x53 ;
  assign n205 = n204 ^ x53 ;
  assign n227 = x47 & ~x48 ;
  assign n228 = ~n205 & n227 ;
  assign n229 = n203 & n228 ;
  assign n230 = n226 & n229 ;
  assign n208 = ~n203 & ~n205 ;
  assign n206 = ~x48 & ~n205 ;
  assign n207 = n203 & n206 ;
  assign n209 = n208 ^ n207 ;
  assign n231 = n230 ^ n209 ;
  assign n232 = x36 & x37 ;
  assign n233 = x38 & x41 ;
  assign n234 = n232 & n233 ;
  assign n235 = x32 & x33 ;
  assign n236 = x34 & x35 ;
  assign n237 = n235 & n236 ;
  assign n238 = n234 & n237 ;
  assign n239 = x57 & x58 ;
  assign n240 = x59 & n239 ;
  assign n241 = x46 & x47 ;
  assign n242 = n241 ^ x47 ;
  assign n243 = x50 & x56 ;
  assign n244 = n243 ^ x50 ;
  assign n245 = n242 & n244 ;
  assign n246 = n240 & n245 ;
  assign n247 = n238 & n246 ;
  assign n254 = n216 & n220 ;
  assign n255 = n254 ^ n220 ;
  assign n256 = n255 ^ x44 ;
  assign n260 = x54 & x55 ;
  assign n261 = x30 & x31 ;
  assign n262 = n260 & n261 ;
  assign n263 = x48 & x49 ;
  assign n264 = n263 ^ x48 ;
  assign n265 = n264 ^ x49 ;
  assign n266 = n212 & n265 ;
  assign n267 = n266 ^ n212 ;
  assign n268 = n267 ^ n212 ;
  assign n269 = n268 ^ n265 ;
  assign n270 = n262 & n269 ;
  assign n271 = n256 & n270 ;
  assign n272 = n271 ^ n270 ;
  assign n277 = n247 & n272 ;
  assign n257 = n256 ^ x45 ;
  assign n248 = n212 & n213 ;
  assign n249 = x44 & x45 ;
  assign n250 = n249 ^ x45 ;
  assign n251 = x43 & n250 ;
  assign n252 = n248 & n251 ;
  assign n253 = n252 ^ n250 ;
  assign n258 = n257 ^ n253 ;
  assign n278 = n226 & n227 ;
  assign n279 = n278 ^ x48 ;
  assign n280 = n258 & n279 ;
  assign n281 = n280 ^ n258 ;
  assign n282 = n277 & n281 ;
  assign n259 = n247 & n258 ;
  assign n273 = x47 & ~x49 ;
  assign n274 = n226 & n273 ;
  assign n275 = n272 & n274 ;
  assign n276 = n259 & n275 ;
  assign n283 = n282 ^ n276 ;
  assign n284 = n231 & n283 ;
  assign n285 = n284 ^ n283 ;
  assign n286 = x52 & ~x53 ;
  assign n287 = n203 & ~n286 ;
  assign n288 = n279 & n287 ;
  assign n289 = x53 & n260 ;
  assign n314 = ~x56 & x59 ;
  assign n315 = n239 & n314 ;
  assign n321 = ~n289 & n315 ;
  assign n297 = x50 ^ x49 ;
  assign n290 = x51 & x52 ;
  assign n291 = n290 ^ x51 ;
  assign n292 = n291 ^ x52 ;
  assign n298 = n297 ^ n292 ;
  assign n299 = n292 ^ x49 ;
  assign n300 = n298 & n299 ;
  assign n301 = n300 ^ n298 ;
  assign n302 = n301 ^ n299 ;
  assign n303 = n302 ^ x50 ;
  assign n296 = n289 ^ x49 ;
  assign n304 = n303 ^ n296 ;
  assign n308 = n227 & ~n304 ;
  assign n309 = n226 & n308 ;
  assign n306 = ~x48 & ~n304 ;
  assign n305 = ~x49 & ~n304 ;
  assign n307 = n306 ^ n305 ;
  assign n310 = n309 ^ n307 ;
  assign n293 = n292 ^ n289 ;
  assign n294 = n289 & n293 ;
  assign n295 = n294 ^ n289 ;
  assign n311 = n310 ^ n295 ;
  assign n312 = n311 ^ n302 ;
  assign n313 = n312 ^ n298 ;
  assign n316 = n295 ^ n289 ;
  assign n317 = n315 & n316 ;
  assign n318 = ~n313 & n317 ;
  assign n319 = n318 ^ n317 ;
  assign n320 = n319 ^ n317 ;
  assign n322 = n321 ^ n320 ;
  assign n323 = n322 ^ n240 ;
  assign n382 = ~x0 & ~x51 ;
  assign n383 = n323 & n382 ;
  assign n384 = n383 ^ n323 ;
  assign n385 = n384 ^ n382 ;
  assign n386 = n288 & n385 ;
  assign n387 = n386 ^ n385 ;
  assign n388 = n285 & n387 ;
  assign n324 = n288 & n323 ;
  assign n325 = n324 ^ n323 ;
  assign n379 = n285 & n325 ;
  assign n380 = n379 ^ n323 ;
  assign n326 = n203 & n205 ;
  assign n327 = x47 & x48 ;
  assign n328 = n326 & n327 ;
  assign n329 = n328 ^ n326 ;
  assign n330 = x33 & x34 ;
  assign n331 = n330 ^ x33 ;
  assign n332 = n331 ^ x34 ;
  assign n333 = x35 & x36 ;
  assign n334 = n333 ^ x35 ;
  assign n335 = n334 ^ x36 ;
  assign n336 = ~n332 & ~n335 ;
  assign n337 = x31 & x32 ;
  assign n338 = n337 ^ x31 ;
  assign n339 = n338 ^ x32 ;
  assign n340 = n260 & ~n339 ;
  assign n341 = n336 & n340 ;
  assign n342 = n329 & n341 ;
  assign n343 = x41 & x43 ;
  assign n344 = n343 ^ x41 ;
  assign n345 = n249 & n344 ;
  assign n346 = x37 & x38 ;
  assign n347 = n346 ^ x37 ;
  assign n348 = n347 ^ x38 ;
  assign n349 = n211 & ~n348 ;
  assign n350 = n345 & n349 ;
  assign n351 = x56 & x57 ;
  assign n352 = n351 ^ x57 ;
  assign n353 = x46 & x51 ;
  assign n354 = n353 ^ x46 ;
  assign n355 = n354 ^ x51 ;
  assign n356 = n352 & ~n355 ;
  assign n357 = x41 & n212 ;
  assign n358 = n357 ^ x41 ;
  assign n359 = n358 ^ x41 ;
  assign n360 = n359 ^ x42 ;
  assign n361 = n356 & n360 ;
  assign n362 = n350 & n361 ;
  assign n363 = n342 & n362 ;
  assign n367 = ~x0 & ~x30 ;
  assign n370 = x48 & n367 ;
  assign n371 = n226 & n370 ;
  assign n372 = n371 ^ n370 ;
  assign n373 = n363 & n372 ;
  assign n364 = x47 & n226 ;
  assign n365 = n364 ^ x47 ;
  assign n366 = n365 ^ x47 ;
  assign n368 = n366 & n367 ;
  assign n369 = n363 & n368 ;
  assign n374 = n373 ^ n369 ;
  assign n377 = n323 & n374 ;
  assign n375 = n325 & n374 ;
  assign n376 = n285 & n375 ;
  assign n378 = n377 ^ n376 ;
  assign n381 = n380 ^ n378 ;
  assign n389 = n388 ^ n381 ;
  assign n414 = n413 ^ n389 ;
  assign n397 = n141 ^ n137 ;
  assign n390 = n137 ^ n110 ;
  assign n391 = ~n137 & n141 ;
  assign n392 = n391 ^ n141 ;
  assign n393 = n392 ^ n110 ;
  assign n394 = n390 & n393 ;
  assign n395 = n394 ^ n390 ;
  assign n396 = n395 ^ n391 ;
  assign n398 = n397 ^ n396 ;
  assign n415 = n414 ^ n398 ;
  assign n419 = n414 ^ n413 ;
  assign n420 = n415 & n419 ;
  assign n421 = n420 ^ n415 ;
  assign n422 = n421 ^ n419 ;
  assign n423 = n422 ^ n414 ;
  assign n424 = n135 & n423 ;
  assign n425 = n424 ^ n135 ;
  assign n426 = n425 ^ n135 ;
  assign n427 = n426 ^ n423 ;
  assign n416 = n415 ^ n413 ;
  assign n417 = n389 & n416 ;
  assign n418 = n417 ^ n416 ;
  assign n428 = n427 ^ n418 ;
  assign n429 = n428 ^ n389 ;
  assign n430 = n429 ^ n135 ;
  assign n431 = n430 ^ n389 ;
  assign n432 = x0 & x30 ;
  assign n433 = x48 & ~n226 ;
  assign n434 = ~n366 & ~n433 ;
  assign n435 = n363 & ~n434 ;
  assign n436 = ~n432 & n435 ;
  assign n437 = n323 & ~n436 ;
  assign n438 = n202 & n437 ;
  assign y0 = ~n202 ;
  assign y1 = ~n431 ;
  assign y2 = n438 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
