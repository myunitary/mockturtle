module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 ;
  assign n33 = ~x24 & ~x25 ;
  assign n34 = ~x26 & ~x27 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x20 & ~x21 ;
  assign n37 = ~x22 & ~x23 ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = x8 & x9 ;
  assign n41 = n40 ^ x8 ;
  assign n42 = n41 ^ x9 ;
  assign n43 = x10 & x11 ;
  assign n44 = n43 ^ x10 ;
  assign n45 = n44 ^ x11 ;
  assign n46 = n42 & n45 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = ~x28 & ~x29 ;
  assign n50 = ~x30 & ~x31 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~n48 & n51 ;
  assign n53 = n39 & n52 ;
  assign n54 = x0 & x1 ;
  assign n55 = n54 ^ x0 ;
  assign n56 = n55 ^ x1 ;
  assign n57 = x2 & x3 ;
  assign n58 = n57 ^ x2 ;
  assign n59 = n58 ^ x3 ;
  assign n60 = n56 & n59 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = x4 & x5 ;
  assign n64 = n63 ^ x4 ;
  assign n65 = n64 ^ x5 ;
  assign n66 = x6 & x7 ;
  assign n67 = n66 ^ x6 ;
  assign n68 = n67 ^ x7 ;
  assign n69 = n65 & n68 ;
  assign n70 = n69 ^ n65 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n62 & ~n71 ;
  assign n73 = x12 & x13 ;
  assign n74 = n73 ^ x12 ;
  assign n75 = n74 ^ x13 ;
  assign n76 = ~x14 & ~x15 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = ~x16 & ~x17 ;
  assign n79 = ~x18 & ~x19 ;
  assign n80 = n78 & n79 ;
  assign n81 = n77 & n80 ;
  assign n82 = n72 & n81 ;
  assign n83 = n53 & n82 ;
  assign n106 = x14 & x15 ;
  assign n107 = n106 ^ x15 ;
  assign n108 = n107 ^ x14 ;
  assign n109 = n75 & n108 ;
  assign n110 = n109 ^ n108 ;
  assign n104 = ~x12 & x13 ;
  assign n105 = n104 ^ x12 ;
  assign n111 = n110 ^ n105 ;
  assign n112 = ~n48 & n111 ;
  assign n100 = ~x10 & x11 ;
  assign n101 = n100 ^ x10 ;
  assign n102 = ~n42 & n101 ;
  assign n98 = ~x8 & x9 ;
  assign n99 = n98 ^ x8 ;
  assign n103 = n102 ^ n99 ;
  assign n113 = n112 ^ n103 ;
  assign n114 = n72 & n113 ;
  assign n92 = ~x6 & x7 ;
  assign n93 = n92 ^ x6 ;
  assign n94 = ~n65 & n93 ;
  assign n90 = ~x4 & x5 ;
  assign n91 = n90 ^ x4 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = ~n62 & n95 ;
  assign n86 = ~x2 & x3 ;
  assign n87 = n86 ^ x2 ;
  assign n88 = ~n56 & n87 ;
  assign n84 = ~x0 & x1 ;
  assign n85 = n84 ^ x0 ;
  assign n89 = n88 ^ n85 ;
  assign n97 = n96 ^ n89 ;
  assign n115 = n114 ^ n97 ;
  assign n164 = n66 & n115 ;
  assign n162 = x22 & x23 ;
  assign n163 = ~n115 & n162 ;
  assign n165 = n164 ^ n163 ;
  assign n160 = x7 & n115 ;
  assign n158 = x23 & n115 ;
  assign n159 = n158 ^ x23 ;
  assign n161 = n160 ^ n159 ;
  assign n166 = n165 ^ n161 ;
  assign n156 = x6 & n115 ;
  assign n154 = x22 & n115 ;
  assign n155 = n154 ^ x22 ;
  assign n157 = n156 ^ n155 ;
  assign n167 = n166 ^ n157 ;
  assign n170 = n63 & n115 ;
  assign n168 = x20 & x21 ;
  assign n169 = ~n115 & n168 ;
  assign n171 = n170 ^ n169 ;
  assign n146 = x5 & n115 ;
  assign n144 = x21 & n115 ;
  assign n145 = n144 ^ x21 ;
  assign n147 = n146 ^ n145 ;
  assign n172 = n171 ^ n147 ;
  assign n150 = x4 & n115 ;
  assign n148 = x20 & n115 ;
  assign n149 = n148 ^ x20 ;
  assign n151 = n150 ^ n149 ;
  assign n173 = n172 ^ n151 ;
  assign n174 = n167 & n173 ;
  assign n175 = n174 ^ n167 ;
  assign n152 = n147 & ~n151 ;
  assign n153 = n152 ^ n151 ;
  assign n176 = n175 ^ n153 ;
  assign n128 = n54 & n115 ;
  assign n126 = x16 & x17 ;
  assign n127 = ~n115 & n126 ;
  assign n129 = n128 ^ n127 ;
  assign n118 = x0 & n115 ;
  assign n116 = x16 & n115 ;
  assign n117 = n116 ^ x16 ;
  assign n119 = n118 ^ n117 ;
  assign n130 = n129 ^ n119 ;
  assign n122 = x1 & n115 ;
  assign n120 = x17 & n115 ;
  assign n121 = n120 ^ x17 ;
  assign n123 = n122 ^ n121 ;
  assign n131 = n130 ^ n123 ;
  assign n179 = n57 & n115 ;
  assign n177 = x18 & x19 ;
  assign n178 = ~n115 & n177 ;
  assign n180 = n179 ^ n178 ;
  assign n134 = x3 & n115 ;
  assign n132 = x19 & n115 ;
  assign n133 = n132 ^ x19 ;
  assign n135 = n134 ^ n133 ;
  assign n181 = n180 ^ n135 ;
  assign n138 = x2 & n115 ;
  assign n136 = x18 & n115 ;
  assign n137 = n136 ^ x18 ;
  assign n139 = n138 ^ n137 ;
  assign n182 = n181 ^ n139 ;
  assign n183 = n131 & n182 ;
  assign n184 = n183 ^ n131 ;
  assign n185 = n184 ^ n182 ;
  assign n186 = n176 & ~n185 ;
  assign n140 = n135 & ~n139 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = ~n131 & n141 ;
  assign n124 = ~n119 & n123 ;
  assign n125 = n124 ^ n119 ;
  assign n143 = n142 ^ n125 ;
  assign n187 = n186 ^ n143 ;
  assign n203 = x10 & n115 ;
  assign n202 = x26 & ~n115 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = n187 & n204 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n206 ^ n139 ;
  assign n209 = x11 & n115 ;
  assign n208 = x27 & ~n115 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n187 & n210 ;
  assign n212 = n211 ^ n210 ;
  assign n213 = n212 ^ n135 ;
  assign n214 = n207 & n213 ;
  assign n215 = n214 ^ n207 ;
  assign n216 = n215 ^ n213 ;
  assign n189 = x8 & n115 ;
  assign n188 = x24 & ~n115 ;
  assign n190 = n189 ^ n188 ;
  assign n191 = n187 & n190 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = n192 ^ n119 ;
  assign n195 = x9 & n115 ;
  assign n194 = x25 & ~n115 ;
  assign n196 = n195 ^ n194 ;
  assign n197 = n187 & n196 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = n198 ^ n123 ;
  assign n217 = n193 & n199 ;
  assign n218 = n217 ^ n193 ;
  assign n219 = n218 ^ n199 ;
  assign n220 = ~n216 & ~n219 ;
  assign n221 = n220 ^ n219 ;
  assign n200 = ~n193 & n199 ;
  assign n201 = n200 ^ n193 ;
  assign n222 = n221 ^ n201 ;
  assign n227 = n147 & n187 ;
  assign n224 = x13 & n115 ;
  assign n223 = x29 & ~n115 ;
  assign n225 = n224 ^ n223 ;
  assign n226 = ~n187 & n225 ;
  assign n228 = n227 ^ n226 ;
  assign n231 = n228 ^ n199 ;
  assign n232 = n231 ^ n228 ;
  assign n233 = ~n193 & ~n232 ;
  assign n229 = n228 ^ n221 ;
  assign n230 = n229 ^ n228 ;
  assign n234 = n233 ^ n230 ;
  assign n239 = n151 & n187 ;
  assign n236 = x12 & n115 ;
  assign n235 = x28 & ~n115 ;
  assign n237 = n236 ^ n235 ;
  assign n238 = ~n187 & n237 ;
  assign n240 = n239 ^ n238 ;
  assign n241 = n240 ^ n193 ;
  assign n242 = ~n228 & ~n241 ;
  assign n243 = n242 ^ n230 ;
  assign n244 = ~n234 & ~n243 ;
  assign n245 = n244 ^ n230 ;
  assign n253 = n157 & n187 ;
  assign n250 = x14 & n115 ;
  assign n249 = x30 & ~n115 ;
  assign n251 = n250 ^ n249 ;
  assign n252 = ~n187 & n251 ;
  assign n254 = n253 ^ n252 ;
  assign n255 = n254 ^ n207 ;
  assign n257 = n255 ^ n254 ;
  assign n256 = n255 ^ n222 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n257 ^ n255 ;
  assign n260 = ~n258 & n259 ;
  assign n261 = n260 ^ n257 ;
  assign n262 = ~n245 & n261 ;
  assign n246 = ~n222 & n240 ;
  assign n247 = n246 ^ n240 ;
  assign n248 = n247 ^ n193 ;
  assign n263 = n262 ^ n248 ;
  assign y0 = 1'b0 ;
  assign y1 = 1'b0 ;
  assign y2 = 1'b0 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = n83 ;
  assign y27 = ~n115 ;
  assign y28 = ~n187 ;
  assign y29 = n222 ;
  assign y30 = ~n245 ;
  assign y31 = ~n263 ;
endmodule
