// Benchmark "bar" written by ABC on Wed Dec 27 23:19:07 2023

module top ( 
    a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15,
    a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29,
    a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43,
    a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57,
    a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71,
    a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85,
    a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99,
    a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111,
    a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123,
    a124, a125, a126, a127, shift0, shift1, shift2, shift3, shift4, shift5,
    shift6,
    ores0, ores1, ores2, ores3, ores4, ores5, ores6, ores7, ores8, ores9,
    ores10, ores11, ores12, ores13, ores14, ores15, ores16, ores17, ores18,
    ores19, ores20, ores21, ores22, ores23, ores24, ores25, ores26, ores27,
    ores28, ores29, ores30, ores31, ores32, ores33, ores34, ores35, ores36,
    ores37, ores38, ores39, ores40, ores41, ores42, ores43, ores44, ores45,
    ores46, ores47, ores48, ores49, ores50, ores51, ores52, ores53, ores54,
    ores55, ores56, ores57, ores58, ores59, ores60, ores61, ores62, ores63,
    ores64, ores65, ores66, ores67, ores68, ores69, ores70, ores71, ores72,
    ores73, ores74, ores75, ores76, ores77, ores78, ores79, ores80, ores81,
    ores82, ores83, ores84, ores85, ores86, ores87, ores88, ores89, ores90,
    ores91, ores92, ores93, ores94, ores95, ores96, ores97, ores98, ores99,
    ores100, ores101, ores102, ores103, ores104, ores105, ores106, ores107,
    ores108, ores109, ores110, ores111, ores112, ores113, ores114, ores115,
    ores116, ores117, ores118, ores119, ores120, ores121, ores122, ores123,
    ores124, ores125, ores126, ores127  );
  input  a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14,
    a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28,
    a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42,
    a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56,
    a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70,
    a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84,
    a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98,
    a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110,
    a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122,
    a123, a124, a125, a126, a127, shift0, shift1, shift2, shift3, shift4,
    shift5, shift6;
  output ores0, ores1, ores2, ores3, ores4, ores5, ores6, ores7, ores8, ores9,
    ores10, ores11, ores12, ores13, ores14, ores15, ores16, ores17, ores18,
    ores19, ores20, ores21, ores22, ores23, ores24, ores25, ores26, ores27,
    ores28, ores29, ores30, ores31, ores32, ores33, ores34, ores35, ores36,
    ores37, ores38, ores39, ores40, ores41, ores42, ores43, ores44, ores45,
    ores46, ores47, ores48, ores49, ores50, ores51, ores52, ores53, ores54,
    ores55, ores56, ores57, ores58, ores59, ores60, ores61, ores62, ores63,
    ores64, ores65, ores66, ores67, ores68, ores69, ores70, ores71, ores72,
    ores73, ores74, ores75, ores76, ores77, ores78, ores79, ores80, ores81,
    ores82, ores83, ores84, ores85, ores86, ores87, ores88, ores89, ores90,
    ores91, ores92, ores93, ores94, ores95, ores96, ores97, ores98, ores99,
    ores100, ores101, ores102, ores103, ores104, ores105, ores106, ores107,
    ores108, ores109, ores110, ores111, ores112, ores113, ores114, ores115,
    ores116, ores117, ores118, ores119, ores120, ores121, ores122, ores123,
    ores124, ores125, ores126, ores127;
  wire new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_,
    new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_,
    new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_,
    new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_,
    new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_,
    new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_,
    new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_,
    new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_,
    new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_,
    new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_,
    new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_,
    new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_,
    new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_,
    new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_,
    new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_,
    new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_,
    new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_,
    new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_,
    new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_,
    new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_,
    new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_,
    new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_,
    new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_,
    new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_,
    new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_,
    new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4540_,
    new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_,
    new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_,
    new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_,
    new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_,
    new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4780_, new_n4781_, new_n4782_,
    new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_,
    new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_,
    new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_,
    new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_,
    new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4960_, new_n4961_, new_n4962_,
    new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_,
    new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_,
    new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_,
    new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_,
    new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_,
    new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5140_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_,
    new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_,
    new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_,
    new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_,
    new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_,
    new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_,
    new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_,
    new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_,
    new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_,
    new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5812_,
    new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5848_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5860_, new_n5861_, new_n5862_,
    new_n5863_, new_n5864_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5884_,
    new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5896_, new_n5897_, new_n5898_,
    new_n5899_, new_n5900_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5956_,
    new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_;
  assign new_n264_ = ~shift6;
  assign new_n265_ = ~shift2;
  assign new_n266_ = ~shift3;
  assign new_n267_ = new_n266_ & new_n265_;
  assign new_n268_ = ~a78;
  assign new_n269_ = ~shift0;
  assign new_n270_ = new_n269_ & new_n268_;
  assign new_n271_ = ~new_n270_;
  assign new_n272_ = ~a77;
  assign new_n273_ = shift0 & new_n272_;
  assign new_n274_ = ~new_n273_;
  assign new_n275_ = new_n274_ & new_n271_;
  assign new_n276_ = ~new_n275_;
  assign new_n277_ = new_n276_ & shift1;
  assign new_n278_ = ~new_n277_;
  assign new_n279_ = ~shift1;
  assign new_n280_ = ~a79;
  assign new_n281_ = shift0 & new_n280_;
  assign new_n282_ = ~new_n281_;
  assign new_n283_ = ~a80;
  assign new_n284_ = new_n269_ & new_n283_;
  assign new_n285_ = ~new_n284_;
  assign new_n286_ = new_n285_ & new_n282_;
  assign new_n287_ = ~new_n286_;
  assign new_n288_ = new_n287_ & new_n279_;
  assign new_n289_ = ~new_n288_;
  assign new_n290_ = new_n289_ & new_n278_;
  assign new_n291_ = new_n290_ & new_n267_;
  assign new_n292_ = ~new_n291_;
  assign new_n293_ = new_n266_ & shift2;
  assign new_n294_ = ~a74;
  assign new_n295_ = new_n269_ & new_n294_;
  assign new_n296_ = ~new_n295_;
  assign new_n297_ = ~a73;
  assign new_n298_ = shift0 & new_n297_;
  assign new_n299_ = ~new_n298_;
  assign new_n300_ = new_n299_ & new_n296_;
  assign new_n301_ = ~new_n300_;
  assign new_n302_ = new_n301_ & shift1;
  assign new_n303_ = ~new_n302_;
  assign new_n304_ = ~a75;
  assign new_n305_ = shift0 & new_n304_;
  assign new_n306_ = ~new_n305_;
  assign new_n307_ = ~a76;
  assign new_n308_ = new_n269_ & new_n307_;
  assign new_n309_ = ~new_n308_;
  assign new_n310_ = new_n309_ & new_n306_;
  assign new_n311_ = ~new_n310_;
  assign new_n312_ = new_n311_ & new_n279_;
  assign new_n313_ = ~new_n312_;
  assign new_n314_ = new_n313_ & new_n303_;
  assign new_n315_ = new_n314_ & new_n293_;
  assign new_n316_ = ~new_n315_;
  assign new_n317_ = new_n316_ & new_n292_;
  assign new_n318_ = shift3 & shift2;
  assign new_n319_ = ~a66;
  assign new_n320_ = new_n269_ & new_n319_;
  assign new_n321_ = ~new_n320_;
  assign new_n322_ = ~a65;
  assign new_n323_ = shift0 & new_n322_;
  assign new_n324_ = ~new_n323_;
  assign new_n325_ = new_n324_ & new_n321_;
  assign new_n326_ = ~new_n325_;
  assign new_n327_ = new_n326_ & shift1;
  assign new_n328_ = ~new_n327_;
  assign new_n329_ = ~a67;
  assign new_n330_ = shift0 & new_n329_;
  assign new_n331_ = ~new_n330_;
  assign new_n332_ = ~a68;
  assign new_n333_ = new_n269_ & new_n332_;
  assign new_n334_ = ~new_n333_;
  assign new_n335_ = new_n334_ & new_n331_;
  assign new_n336_ = ~new_n335_;
  assign new_n337_ = new_n336_ & new_n279_;
  assign new_n338_ = ~new_n337_;
  assign new_n339_ = new_n338_ & new_n328_;
  assign new_n340_ = new_n339_ & new_n318_;
  assign new_n341_ = ~new_n340_;
  assign new_n342_ = shift3 & new_n265_;
  assign new_n343_ = ~a70;
  assign new_n344_ = new_n269_ & new_n343_;
  assign new_n345_ = ~new_n344_;
  assign new_n346_ = ~a69;
  assign new_n347_ = shift0 & new_n346_;
  assign new_n348_ = ~new_n347_;
  assign new_n349_ = new_n348_ & new_n345_;
  assign new_n350_ = ~new_n349_;
  assign new_n351_ = new_n350_ & shift1;
  assign new_n352_ = ~new_n351_;
  assign new_n353_ = ~a71;
  assign new_n354_ = shift0 & new_n353_;
  assign new_n355_ = ~new_n354_;
  assign new_n356_ = ~a72;
  assign new_n357_ = new_n269_ & new_n356_;
  assign new_n358_ = ~new_n357_;
  assign new_n359_ = new_n358_ & new_n355_;
  assign new_n360_ = ~new_n359_;
  assign new_n361_ = new_n360_ & new_n279_;
  assign new_n362_ = ~new_n361_;
  assign new_n363_ = new_n362_ & new_n352_;
  assign new_n364_ = new_n363_ & new_n342_;
  assign new_n365_ = ~new_n364_;
  assign new_n366_ = new_n365_ & new_n341_;
  assign new_n367_ = new_n366_ & new_n317_;
  assign new_n368_ = ~new_n367_;
  assign new_n369_ = shift5 & shift4;
  assign new_n370_ = new_n369_ & new_n368_;
  assign new_n371_ = ~new_n370_;
  assign new_n372_ = ~a94;
  assign new_n373_ = new_n269_ & new_n372_;
  assign new_n374_ = ~new_n373_;
  assign new_n375_ = ~a93;
  assign new_n376_ = shift0 & new_n375_;
  assign new_n377_ = ~new_n376_;
  assign new_n378_ = new_n377_ & new_n374_;
  assign new_n379_ = ~new_n378_;
  assign new_n380_ = new_n379_ & shift1;
  assign new_n381_ = ~new_n380_;
  assign new_n382_ = ~a95;
  assign new_n383_ = shift0 & new_n382_;
  assign new_n384_ = ~new_n383_;
  assign new_n385_ = ~a96;
  assign new_n386_ = new_n269_ & new_n385_;
  assign new_n387_ = ~new_n386_;
  assign new_n388_ = new_n387_ & new_n384_;
  assign new_n389_ = ~new_n388_;
  assign new_n390_ = new_n389_ & new_n279_;
  assign new_n391_ = ~new_n390_;
  assign new_n392_ = new_n391_ & new_n381_;
  assign new_n393_ = new_n392_ & new_n267_;
  assign new_n394_ = ~new_n393_;
  assign new_n395_ = ~a90;
  assign new_n396_ = new_n269_ & new_n395_;
  assign new_n397_ = ~new_n396_;
  assign new_n398_ = ~a89;
  assign new_n399_ = shift0 & new_n398_;
  assign new_n400_ = ~new_n399_;
  assign new_n401_ = new_n400_ & new_n397_;
  assign new_n402_ = ~new_n401_;
  assign new_n403_ = new_n402_ & shift1;
  assign new_n404_ = ~new_n403_;
  assign new_n405_ = ~a91;
  assign new_n406_ = shift0 & new_n405_;
  assign new_n407_ = ~new_n406_;
  assign new_n408_ = ~a92;
  assign new_n409_ = new_n269_ & new_n408_;
  assign new_n410_ = ~new_n409_;
  assign new_n411_ = new_n410_ & new_n407_;
  assign new_n412_ = ~new_n411_;
  assign new_n413_ = new_n412_ & new_n279_;
  assign new_n414_ = ~new_n413_;
  assign new_n415_ = new_n414_ & new_n404_;
  assign new_n416_ = new_n415_ & new_n293_;
  assign new_n417_ = ~new_n416_;
  assign new_n418_ = new_n417_ & new_n394_;
  assign new_n419_ = ~a82;
  assign new_n420_ = new_n269_ & new_n419_;
  assign new_n421_ = ~new_n420_;
  assign new_n422_ = ~a81;
  assign new_n423_ = shift0 & new_n422_;
  assign new_n424_ = ~new_n423_;
  assign new_n425_ = new_n424_ & new_n421_;
  assign new_n426_ = ~new_n425_;
  assign new_n427_ = new_n426_ & shift1;
  assign new_n428_ = ~new_n427_;
  assign new_n429_ = ~a83;
  assign new_n430_ = shift0 & new_n429_;
  assign new_n431_ = ~new_n430_;
  assign new_n432_ = ~a84;
  assign new_n433_ = new_n269_ & new_n432_;
  assign new_n434_ = ~new_n433_;
  assign new_n435_ = new_n434_ & new_n431_;
  assign new_n436_ = ~new_n435_;
  assign new_n437_ = new_n436_ & new_n279_;
  assign new_n438_ = ~new_n437_;
  assign new_n439_ = new_n438_ & new_n428_;
  assign new_n440_ = new_n439_ & new_n318_;
  assign new_n441_ = ~new_n440_;
  assign new_n442_ = ~a86;
  assign new_n443_ = new_n269_ & new_n442_;
  assign new_n444_ = ~new_n443_;
  assign new_n445_ = ~a85;
  assign new_n446_ = shift0 & new_n445_;
  assign new_n447_ = ~new_n446_;
  assign new_n448_ = new_n447_ & new_n444_;
  assign new_n449_ = ~new_n448_;
  assign new_n450_ = new_n449_ & shift1;
  assign new_n451_ = ~new_n450_;
  assign new_n452_ = ~a87;
  assign new_n453_ = shift0 & new_n452_;
  assign new_n454_ = ~new_n453_;
  assign new_n455_ = ~a88;
  assign new_n456_ = new_n269_ & new_n455_;
  assign new_n457_ = ~new_n456_;
  assign new_n458_ = new_n457_ & new_n454_;
  assign new_n459_ = ~new_n458_;
  assign new_n460_ = new_n459_ & new_n279_;
  assign new_n461_ = ~new_n460_;
  assign new_n462_ = new_n461_ & new_n451_;
  assign new_n463_ = new_n462_ & new_n342_;
  assign new_n464_ = ~new_n463_;
  assign new_n465_ = new_n464_ & new_n441_;
  assign new_n466_ = new_n465_ & new_n418_;
  assign new_n467_ = ~new_n466_;
  assign new_n468_ = ~shift4;
  assign new_n469_ = shift5 & new_n468_;
  assign new_n470_ = new_n469_ & new_n467_;
  assign new_n471_ = ~new_n470_;
  assign new_n472_ = new_n471_ & new_n371_;
  assign new_n473_ = ~a126;
  assign new_n474_ = new_n269_ & new_n473_;
  assign new_n475_ = ~new_n474_;
  assign new_n476_ = ~a125;
  assign new_n477_ = shift0 & new_n476_;
  assign new_n478_ = ~new_n477_;
  assign new_n479_ = new_n478_ & new_n475_;
  assign new_n480_ = ~new_n479_;
  assign new_n481_ = new_n480_ & shift1;
  assign new_n482_ = ~new_n481_;
  assign new_n483_ = ~a127;
  assign new_n484_ = shift0 & new_n483_;
  assign new_n485_ = ~new_n484_;
  assign new_n486_ = ~a0;
  assign new_n487_ = new_n269_ & new_n486_;
  assign new_n488_ = ~new_n487_;
  assign new_n489_ = new_n488_ & new_n485_;
  assign new_n490_ = ~new_n489_;
  assign new_n491_ = new_n490_ & new_n279_;
  assign new_n492_ = ~new_n491_;
  assign new_n493_ = new_n492_ & new_n482_;
  assign new_n494_ = new_n493_ & new_n267_;
  assign new_n495_ = ~new_n494_;
  assign new_n496_ = ~a122;
  assign new_n497_ = new_n269_ & new_n496_;
  assign new_n498_ = ~new_n497_;
  assign new_n499_ = ~a121;
  assign new_n500_ = shift0 & new_n499_;
  assign new_n501_ = ~new_n500_;
  assign new_n502_ = new_n501_ & new_n498_;
  assign new_n503_ = ~new_n502_;
  assign new_n504_ = new_n503_ & shift1;
  assign new_n505_ = ~new_n504_;
  assign new_n506_ = ~a123;
  assign new_n507_ = shift0 & new_n506_;
  assign new_n508_ = ~new_n507_;
  assign new_n509_ = ~a124;
  assign new_n510_ = new_n269_ & new_n509_;
  assign new_n511_ = ~new_n510_;
  assign new_n512_ = new_n511_ & new_n508_;
  assign new_n513_ = ~new_n512_;
  assign new_n514_ = new_n513_ & new_n279_;
  assign new_n515_ = ~new_n514_;
  assign new_n516_ = new_n515_ & new_n505_;
  assign new_n517_ = new_n516_ & new_n293_;
  assign new_n518_ = ~new_n517_;
  assign new_n519_ = new_n518_ & new_n495_;
  assign new_n520_ = ~a114;
  assign new_n521_ = new_n269_ & new_n520_;
  assign new_n522_ = ~new_n521_;
  assign new_n523_ = ~a113;
  assign new_n524_ = shift0 & new_n523_;
  assign new_n525_ = ~new_n524_;
  assign new_n526_ = new_n525_ & new_n522_;
  assign new_n527_ = ~new_n526_;
  assign new_n528_ = new_n527_ & shift1;
  assign new_n529_ = ~new_n528_;
  assign new_n530_ = ~a115;
  assign new_n531_ = shift0 & new_n530_;
  assign new_n532_ = ~new_n531_;
  assign new_n533_ = ~a116;
  assign new_n534_ = new_n269_ & new_n533_;
  assign new_n535_ = ~new_n534_;
  assign new_n536_ = new_n535_ & new_n532_;
  assign new_n537_ = ~new_n536_;
  assign new_n538_ = new_n537_ & new_n279_;
  assign new_n539_ = ~new_n538_;
  assign new_n540_ = new_n539_ & new_n529_;
  assign new_n541_ = new_n540_ & new_n318_;
  assign new_n542_ = ~new_n541_;
  assign new_n543_ = ~a118;
  assign new_n544_ = new_n269_ & new_n543_;
  assign new_n545_ = ~new_n544_;
  assign new_n546_ = ~a117;
  assign new_n547_ = shift0 & new_n546_;
  assign new_n548_ = ~new_n547_;
  assign new_n549_ = new_n548_ & new_n545_;
  assign new_n550_ = ~new_n549_;
  assign new_n551_ = new_n550_ & shift1;
  assign new_n552_ = ~new_n551_;
  assign new_n553_ = ~a119;
  assign new_n554_ = shift0 & new_n553_;
  assign new_n555_ = ~new_n554_;
  assign new_n556_ = ~a120;
  assign new_n557_ = new_n269_ & new_n556_;
  assign new_n558_ = ~new_n557_;
  assign new_n559_ = new_n558_ & new_n555_;
  assign new_n560_ = ~new_n559_;
  assign new_n561_ = new_n560_ & new_n279_;
  assign new_n562_ = ~new_n561_;
  assign new_n563_ = new_n562_ & new_n552_;
  assign new_n564_ = new_n563_ & new_n342_;
  assign new_n565_ = ~new_n564_;
  assign new_n566_ = new_n565_ & new_n542_;
  assign new_n567_ = new_n566_ & new_n519_;
  assign new_n568_ = ~new_n567_;
  assign new_n569_ = ~shift5;
  assign new_n570_ = new_n569_ & new_n468_;
  assign new_n571_ = new_n570_ & new_n568_;
  assign new_n572_ = ~new_n571_;
  assign new_n573_ = ~a110;
  assign new_n574_ = new_n269_ & new_n573_;
  assign new_n575_ = ~new_n574_;
  assign new_n576_ = ~a109;
  assign new_n577_ = shift0 & new_n576_;
  assign new_n578_ = ~new_n577_;
  assign new_n579_ = new_n578_ & new_n575_;
  assign new_n580_ = ~new_n579_;
  assign new_n581_ = new_n580_ & shift1;
  assign new_n582_ = ~new_n581_;
  assign new_n583_ = ~a111;
  assign new_n584_ = shift0 & new_n583_;
  assign new_n585_ = ~new_n584_;
  assign new_n586_ = ~a112;
  assign new_n587_ = new_n269_ & new_n586_;
  assign new_n588_ = ~new_n587_;
  assign new_n589_ = new_n588_ & new_n585_;
  assign new_n590_ = ~new_n589_;
  assign new_n591_ = new_n590_ & new_n279_;
  assign new_n592_ = ~new_n591_;
  assign new_n593_ = new_n592_ & new_n582_;
  assign new_n594_ = new_n593_ & new_n267_;
  assign new_n595_ = ~new_n594_;
  assign new_n596_ = ~a106;
  assign new_n597_ = new_n269_ & new_n596_;
  assign new_n598_ = ~new_n597_;
  assign new_n599_ = ~a105;
  assign new_n600_ = shift0 & new_n599_;
  assign new_n601_ = ~new_n600_;
  assign new_n602_ = new_n601_ & new_n598_;
  assign new_n603_ = ~new_n602_;
  assign new_n604_ = new_n603_ & shift1;
  assign new_n605_ = ~new_n604_;
  assign new_n606_ = ~a107;
  assign new_n607_ = shift0 & new_n606_;
  assign new_n608_ = ~new_n607_;
  assign new_n609_ = ~a108;
  assign new_n610_ = new_n269_ & new_n609_;
  assign new_n611_ = ~new_n610_;
  assign new_n612_ = new_n611_ & new_n608_;
  assign new_n613_ = ~new_n612_;
  assign new_n614_ = new_n613_ & new_n279_;
  assign new_n615_ = ~new_n614_;
  assign new_n616_ = new_n615_ & new_n605_;
  assign new_n617_ = new_n616_ & new_n293_;
  assign new_n618_ = ~new_n617_;
  assign new_n619_ = new_n618_ & new_n595_;
  assign new_n620_ = ~a98;
  assign new_n621_ = new_n269_ & new_n620_;
  assign new_n622_ = ~new_n621_;
  assign new_n623_ = ~a97;
  assign new_n624_ = shift0 & new_n623_;
  assign new_n625_ = ~new_n624_;
  assign new_n626_ = new_n625_ & new_n622_;
  assign new_n627_ = ~new_n626_;
  assign new_n628_ = new_n627_ & shift1;
  assign new_n629_ = ~new_n628_;
  assign new_n630_ = ~a99;
  assign new_n631_ = shift0 & new_n630_;
  assign new_n632_ = ~new_n631_;
  assign new_n633_ = ~a100;
  assign new_n634_ = new_n269_ & new_n633_;
  assign new_n635_ = ~new_n634_;
  assign new_n636_ = new_n635_ & new_n632_;
  assign new_n637_ = ~new_n636_;
  assign new_n638_ = new_n637_ & new_n279_;
  assign new_n639_ = ~new_n638_;
  assign new_n640_ = new_n639_ & new_n629_;
  assign new_n641_ = new_n640_ & new_n318_;
  assign new_n642_ = ~new_n641_;
  assign new_n643_ = ~a102;
  assign new_n644_ = new_n269_ & new_n643_;
  assign new_n645_ = ~new_n644_;
  assign new_n646_ = ~a101;
  assign new_n647_ = shift0 & new_n646_;
  assign new_n648_ = ~new_n647_;
  assign new_n649_ = new_n648_ & new_n645_;
  assign new_n650_ = ~new_n649_;
  assign new_n651_ = new_n650_ & shift1;
  assign new_n652_ = ~new_n651_;
  assign new_n653_ = ~a103;
  assign new_n654_ = shift0 & new_n653_;
  assign new_n655_ = ~new_n654_;
  assign new_n656_ = ~a104;
  assign new_n657_ = new_n269_ & new_n656_;
  assign new_n658_ = ~new_n657_;
  assign new_n659_ = new_n658_ & new_n655_;
  assign new_n660_ = ~new_n659_;
  assign new_n661_ = new_n660_ & new_n279_;
  assign new_n662_ = ~new_n661_;
  assign new_n663_ = new_n662_ & new_n652_;
  assign new_n664_ = new_n663_ & new_n342_;
  assign new_n665_ = ~new_n664_;
  assign new_n666_ = new_n665_ & new_n642_;
  assign new_n667_ = new_n666_ & new_n619_;
  assign new_n668_ = ~new_n667_;
  assign new_n669_ = new_n569_ & shift4;
  assign new_n670_ = new_n669_ & new_n668_;
  assign new_n671_ = ~new_n670_;
  assign new_n672_ = new_n671_ & new_n572_;
  assign new_n673_ = new_n672_ & new_n472_;
  assign new_n674_ = ~new_n673_;
  assign new_n675_ = new_n674_ & new_n264_;
  assign new_n676_ = ~new_n675_;
  assign new_n677_ = ~a14;
  assign new_n678_ = new_n269_ & new_n677_;
  assign new_n679_ = ~new_n678_;
  assign new_n680_ = ~a13;
  assign new_n681_ = shift0 & new_n680_;
  assign new_n682_ = ~new_n681_;
  assign new_n683_ = new_n682_ & new_n679_;
  assign new_n684_ = ~new_n683_;
  assign new_n685_ = new_n684_ & shift1;
  assign new_n686_ = ~new_n685_;
  assign new_n687_ = ~a15;
  assign new_n688_ = shift0 & new_n687_;
  assign new_n689_ = ~new_n688_;
  assign new_n690_ = ~a16;
  assign new_n691_ = new_n269_ & new_n690_;
  assign new_n692_ = ~new_n691_;
  assign new_n693_ = new_n692_ & new_n689_;
  assign new_n694_ = ~new_n693_;
  assign new_n695_ = new_n694_ & new_n279_;
  assign new_n696_ = ~new_n695_;
  assign new_n697_ = new_n696_ & new_n686_;
  assign new_n698_ = new_n697_ & new_n267_;
  assign new_n699_ = ~new_n698_;
  assign new_n700_ = ~a10;
  assign new_n701_ = new_n269_ & new_n700_;
  assign new_n702_ = ~new_n701_;
  assign new_n703_ = ~a9;
  assign new_n704_ = shift0 & new_n703_;
  assign new_n705_ = ~new_n704_;
  assign new_n706_ = new_n705_ & new_n702_;
  assign new_n707_ = ~new_n706_;
  assign new_n708_ = new_n707_ & shift1;
  assign new_n709_ = ~new_n708_;
  assign new_n710_ = ~a11;
  assign new_n711_ = shift0 & new_n710_;
  assign new_n712_ = ~new_n711_;
  assign new_n713_ = ~a12;
  assign new_n714_ = new_n269_ & new_n713_;
  assign new_n715_ = ~new_n714_;
  assign new_n716_ = new_n715_ & new_n712_;
  assign new_n717_ = ~new_n716_;
  assign new_n718_ = new_n717_ & new_n279_;
  assign new_n719_ = ~new_n718_;
  assign new_n720_ = new_n719_ & new_n709_;
  assign new_n721_ = new_n720_ & new_n293_;
  assign new_n722_ = ~new_n721_;
  assign new_n723_ = new_n722_ & new_n699_;
  assign new_n724_ = ~a2;
  assign new_n725_ = new_n269_ & new_n724_;
  assign new_n726_ = ~new_n725_;
  assign new_n727_ = ~a1;
  assign new_n728_ = shift0 & new_n727_;
  assign new_n729_ = ~new_n728_;
  assign new_n730_ = new_n729_ & new_n726_;
  assign new_n731_ = ~new_n730_;
  assign new_n732_ = new_n731_ & shift1;
  assign new_n733_ = ~new_n732_;
  assign new_n734_ = ~a3;
  assign new_n735_ = shift0 & new_n734_;
  assign new_n736_ = ~new_n735_;
  assign new_n737_ = ~a4;
  assign new_n738_ = new_n269_ & new_n737_;
  assign new_n739_ = ~new_n738_;
  assign new_n740_ = new_n739_ & new_n736_;
  assign new_n741_ = ~new_n740_;
  assign new_n742_ = new_n741_ & new_n279_;
  assign new_n743_ = ~new_n742_;
  assign new_n744_ = new_n743_ & new_n733_;
  assign new_n745_ = new_n744_ & new_n318_;
  assign new_n746_ = ~new_n745_;
  assign new_n747_ = ~a6;
  assign new_n748_ = new_n269_ & new_n747_;
  assign new_n749_ = ~new_n748_;
  assign new_n750_ = ~a5;
  assign new_n751_ = shift0 & new_n750_;
  assign new_n752_ = ~new_n751_;
  assign new_n753_ = new_n752_ & new_n749_;
  assign new_n754_ = ~new_n753_;
  assign new_n755_ = new_n754_ & shift1;
  assign new_n756_ = ~new_n755_;
  assign new_n757_ = ~a7;
  assign new_n758_ = shift0 & new_n757_;
  assign new_n759_ = ~new_n758_;
  assign new_n760_ = ~a8;
  assign new_n761_ = new_n269_ & new_n760_;
  assign new_n762_ = ~new_n761_;
  assign new_n763_ = new_n762_ & new_n759_;
  assign new_n764_ = ~new_n763_;
  assign new_n765_ = new_n764_ & new_n279_;
  assign new_n766_ = ~new_n765_;
  assign new_n767_ = new_n766_ & new_n756_;
  assign new_n768_ = new_n767_ & new_n342_;
  assign new_n769_ = ~new_n768_;
  assign new_n770_ = new_n769_ & new_n746_;
  assign new_n771_ = new_n770_ & new_n723_;
  assign new_n772_ = ~new_n771_;
  assign new_n773_ = new_n772_ & new_n369_;
  assign new_n774_ = ~new_n773_;
  assign new_n775_ = ~a30;
  assign new_n776_ = new_n269_ & new_n775_;
  assign new_n777_ = ~new_n776_;
  assign new_n778_ = ~a29;
  assign new_n779_ = shift0 & new_n778_;
  assign new_n780_ = ~new_n779_;
  assign new_n781_ = new_n780_ & new_n777_;
  assign new_n782_ = ~new_n781_;
  assign new_n783_ = new_n782_ & shift1;
  assign new_n784_ = ~new_n783_;
  assign new_n785_ = ~a31;
  assign new_n786_ = shift0 & new_n785_;
  assign new_n787_ = ~new_n786_;
  assign new_n788_ = ~a32;
  assign new_n789_ = new_n269_ & new_n788_;
  assign new_n790_ = ~new_n789_;
  assign new_n791_ = new_n790_ & new_n787_;
  assign new_n792_ = ~new_n791_;
  assign new_n793_ = new_n792_ & new_n279_;
  assign new_n794_ = ~new_n793_;
  assign new_n795_ = new_n794_ & new_n784_;
  assign new_n796_ = new_n795_ & new_n267_;
  assign new_n797_ = ~new_n796_;
  assign new_n798_ = ~a26;
  assign new_n799_ = new_n269_ & new_n798_;
  assign new_n800_ = ~new_n799_;
  assign new_n801_ = ~a25;
  assign new_n802_ = shift0 & new_n801_;
  assign new_n803_ = ~new_n802_;
  assign new_n804_ = new_n803_ & new_n800_;
  assign new_n805_ = ~new_n804_;
  assign new_n806_ = new_n805_ & shift1;
  assign new_n807_ = ~new_n806_;
  assign new_n808_ = ~a27;
  assign new_n809_ = shift0 & new_n808_;
  assign new_n810_ = ~new_n809_;
  assign new_n811_ = ~a28;
  assign new_n812_ = new_n269_ & new_n811_;
  assign new_n813_ = ~new_n812_;
  assign new_n814_ = new_n813_ & new_n810_;
  assign new_n815_ = ~new_n814_;
  assign new_n816_ = new_n815_ & new_n279_;
  assign new_n817_ = ~new_n816_;
  assign new_n818_ = new_n817_ & new_n807_;
  assign new_n819_ = new_n818_ & new_n293_;
  assign new_n820_ = ~new_n819_;
  assign new_n821_ = new_n820_ & new_n797_;
  assign new_n822_ = ~a18;
  assign new_n823_ = new_n269_ & new_n822_;
  assign new_n824_ = ~new_n823_;
  assign new_n825_ = ~a17;
  assign new_n826_ = shift0 & new_n825_;
  assign new_n827_ = ~new_n826_;
  assign new_n828_ = new_n827_ & new_n824_;
  assign new_n829_ = ~new_n828_;
  assign new_n830_ = new_n829_ & shift1;
  assign new_n831_ = ~new_n830_;
  assign new_n832_ = ~a19;
  assign new_n833_ = shift0 & new_n832_;
  assign new_n834_ = ~new_n833_;
  assign new_n835_ = ~a20;
  assign new_n836_ = new_n269_ & new_n835_;
  assign new_n837_ = ~new_n836_;
  assign new_n838_ = new_n837_ & new_n834_;
  assign new_n839_ = ~new_n838_;
  assign new_n840_ = new_n839_ & new_n279_;
  assign new_n841_ = ~new_n840_;
  assign new_n842_ = new_n841_ & new_n831_;
  assign new_n843_ = new_n842_ & new_n318_;
  assign new_n844_ = ~new_n843_;
  assign new_n845_ = ~a22;
  assign new_n846_ = new_n269_ & new_n845_;
  assign new_n847_ = ~new_n846_;
  assign new_n848_ = ~a21;
  assign new_n849_ = shift0 & new_n848_;
  assign new_n850_ = ~new_n849_;
  assign new_n851_ = new_n850_ & new_n847_;
  assign new_n852_ = ~new_n851_;
  assign new_n853_ = new_n852_ & shift1;
  assign new_n854_ = ~new_n853_;
  assign new_n855_ = ~a23;
  assign new_n856_ = shift0 & new_n855_;
  assign new_n857_ = ~new_n856_;
  assign new_n858_ = ~a24;
  assign new_n859_ = new_n269_ & new_n858_;
  assign new_n860_ = ~new_n859_;
  assign new_n861_ = new_n860_ & new_n857_;
  assign new_n862_ = ~new_n861_;
  assign new_n863_ = new_n862_ & new_n279_;
  assign new_n864_ = ~new_n863_;
  assign new_n865_ = new_n864_ & new_n854_;
  assign new_n866_ = new_n865_ & new_n342_;
  assign new_n867_ = ~new_n866_;
  assign new_n868_ = new_n867_ & new_n844_;
  assign new_n869_ = new_n868_ & new_n821_;
  assign new_n870_ = ~new_n869_;
  assign new_n871_ = new_n870_ & new_n469_;
  assign new_n872_ = ~new_n871_;
  assign new_n873_ = new_n872_ & new_n774_;
  assign new_n874_ = ~a62;
  assign new_n875_ = new_n269_ & new_n874_;
  assign new_n876_ = ~new_n875_;
  assign new_n877_ = ~a61;
  assign new_n878_ = shift0 & new_n877_;
  assign new_n879_ = ~new_n878_;
  assign new_n880_ = new_n879_ & new_n876_;
  assign new_n881_ = ~new_n880_;
  assign new_n882_ = new_n881_ & shift1;
  assign new_n883_ = ~new_n882_;
  assign new_n884_ = ~a63;
  assign new_n885_ = shift0 & new_n884_;
  assign new_n886_ = ~new_n885_;
  assign new_n887_ = ~a64;
  assign new_n888_ = new_n269_ & new_n887_;
  assign new_n889_ = ~new_n888_;
  assign new_n890_ = new_n889_ & new_n886_;
  assign new_n891_ = ~new_n890_;
  assign new_n892_ = new_n891_ & new_n279_;
  assign new_n893_ = ~new_n892_;
  assign new_n894_ = new_n893_ & new_n883_;
  assign new_n895_ = new_n894_ & new_n267_;
  assign new_n896_ = ~new_n895_;
  assign new_n897_ = ~a58;
  assign new_n898_ = new_n269_ & new_n897_;
  assign new_n899_ = ~new_n898_;
  assign new_n900_ = ~a57;
  assign new_n901_ = shift0 & new_n900_;
  assign new_n902_ = ~new_n901_;
  assign new_n903_ = new_n902_ & new_n899_;
  assign new_n904_ = ~new_n903_;
  assign new_n905_ = new_n904_ & shift1;
  assign new_n906_ = ~new_n905_;
  assign new_n907_ = ~a59;
  assign new_n908_ = shift0 & new_n907_;
  assign new_n909_ = ~new_n908_;
  assign new_n910_ = ~a60;
  assign new_n911_ = new_n269_ & new_n910_;
  assign new_n912_ = ~new_n911_;
  assign new_n913_ = new_n912_ & new_n909_;
  assign new_n914_ = ~new_n913_;
  assign new_n915_ = new_n914_ & new_n279_;
  assign new_n916_ = ~new_n915_;
  assign new_n917_ = new_n916_ & new_n906_;
  assign new_n918_ = new_n917_ & new_n293_;
  assign new_n919_ = ~new_n918_;
  assign new_n920_ = new_n919_ & new_n896_;
  assign new_n921_ = ~a50;
  assign new_n922_ = new_n269_ & new_n921_;
  assign new_n923_ = ~new_n922_;
  assign new_n924_ = ~a49;
  assign new_n925_ = shift0 & new_n924_;
  assign new_n926_ = ~new_n925_;
  assign new_n927_ = new_n926_ & new_n923_;
  assign new_n928_ = ~new_n927_;
  assign new_n929_ = new_n928_ & shift1;
  assign new_n930_ = ~new_n929_;
  assign new_n931_ = ~a51;
  assign new_n932_ = shift0 & new_n931_;
  assign new_n933_ = ~new_n932_;
  assign new_n934_ = ~a52;
  assign new_n935_ = new_n269_ & new_n934_;
  assign new_n936_ = ~new_n935_;
  assign new_n937_ = new_n936_ & new_n933_;
  assign new_n938_ = ~new_n937_;
  assign new_n939_ = new_n938_ & new_n279_;
  assign new_n940_ = ~new_n939_;
  assign new_n941_ = new_n940_ & new_n930_;
  assign new_n942_ = new_n941_ & new_n318_;
  assign new_n943_ = ~new_n942_;
  assign new_n944_ = ~a54;
  assign new_n945_ = new_n269_ & new_n944_;
  assign new_n946_ = ~new_n945_;
  assign new_n947_ = ~a53;
  assign new_n948_ = shift0 & new_n947_;
  assign new_n949_ = ~new_n948_;
  assign new_n950_ = new_n949_ & new_n946_;
  assign new_n951_ = ~new_n950_;
  assign new_n952_ = new_n951_ & shift1;
  assign new_n953_ = ~new_n952_;
  assign new_n954_ = ~a55;
  assign new_n955_ = shift0 & new_n954_;
  assign new_n956_ = ~new_n955_;
  assign new_n957_ = ~a56;
  assign new_n958_ = new_n269_ & new_n957_;
  assign new_n959_ = ~new_n958_;
  assign new_n960_ = new_n959_ & new_n956_;
  assign new_n961_ = ~new_n960_;
  assign new_n962_ = new_n961_ & new_n279_;
  assign new_n963_ = ~new_n962_;
  assign new_n964_ = new_n963_ & new_n953_;
  assign new_n965_ = new_n964_ & new_n342_;
  assign new_n966_ = ~new_n965_;
  assign new_n967_ = new_n966_ & new_n943_;
  assign new_n968_ = new_n967_ & new_n920_;
  assign new_n969_ = ~new_n968_;
  assign new_n970_ = new_n969_ & new_n570_;
  assign new_n971_ = ~new_n970_;
  assign new_n972_ = ~a46;
  assign new_n973_ = new_n269_ & new_n972_;
  assign new_n974_ = ~new_n973_;
  assign new_n975_ = ~a45;
  assign new_n976_ = shift0 & new_n975_;
  assign new_n977_ = ~new_n976_;
  assign new_n978_ = new_n977_ & new_n974_;
  assign new_n979_ = ~new_n978_;
  assign new_n980_ = new_n979_ & shift1;
  assign new_n981_ = ~new_n980_;
  assign new_n982_ = ~a47;
  assign new_n983_ = shift0 & new_n982_;
  assign new_n984_ = ~new_n983_;
  assign new_n985_ = ~a48;
  assign new_n986_ = new_n269_ & new_n985_;
  assign new_n987_ = ~new_n986_;
  assign new_n988_ = new_n987_ & new_n984_;
  assign new_n989_ = ~new_n988_;
  assign new_n990_ = new_n989_ & new_n279_;
  assign new_n991_ = ~new_n990_;
  assign new_n992_ = new_n991_ & new_n981_;
  assign new_n993_ = new_n992_ & new_n267_;
  assign new_n994_ = ~new_n993_;
  assign new_n995_ = ~a42;
  assign new_n996_ = new_n269_ & new_n995_;
  assign new_n997_ = ~new_n996_;
  assign new_n998_ = ~a41;
  assign new_n999_ = shift0 & new_n998_;
  assign new_n1000_ = ~new_n999_;
  assign new_n1001_ = new_n1000_ & new_n997_;
  assign new_n1002_ = ~new_n1001_;
  assign new_n1003_ = new_n1002_ & shift1;
  assign new_n1004_ = ~new_n1003_;
  assign new_n1005_ = ~a43;
  assign new_n1006_ = shift0 & new_n1005_;
  assign new_n1007_ = ~new_n1006_;
  assign new_n1008_ = ~a44;
  assign new_n1009_ = new_n269_ & new_n1008_;
  assign new_n1010_ = ~new_n1009_;
  assign new_n1011_ = new_n1010_ & new_n1007_;
  assign new_n1012_ = ~new_n1011_;
  assign new_n1013_ = new_n1012_ & new_n279_;
  assign new_n1014_ = ~new_n1013_;
  assign new_n1015_ = new_n1014_ & new_n1004_;
  assign new_n1016_ = new_n1015_ & new_n293_;
  assign new_n1017_ = ~new_n1016_;
  assign new_n1018_ = new_n1017_ & new_n994_;
  assign new_n1019_ = ~a34;
  assign new_n1020_ = new_n269_ & new_n1019_;
  assign new_n1021_ = ~new_n1020_;
  assign new_n1022_ = ~a33;
  assign new_n1023_ = shift0 & new_n1022_;
  assign new_n1024_ = ~new_n1023_;
  assign new_n1025_ = new_n1024_ & new_n1021_;
  assign new_n1026_ = ~new_n1025_;
  assign new_n1027_ = new_n1026_ & shift1;
  assign new_n1028_ = ~new_n1027_;
  assign new_n1029_ = ~a35;
  assign new_n1030_ = shift0 & new_n1029_;
  assign new_n1031_ = ~new_n1030_;
  assign new_n1032_ = ~a36;
  assign new_n1033_ = new_n269_ & new_n1032_;
  assign new_n1034_ = ~new_n1033_;
  assign new_n1035_ = new_n1034_ & new_n1031_;
  assign new_n1036_ = ~new_n1035_;
  assign new_n1037_ = new_n1036_ & new_n279_;
  assign new_n1038_ = ~new_n1037_;
  assign new_n1039_ = new_n1038_ & new_n1028_;
  assign new_n1040_ = new_n1039_ & new_n318_;
  assign new_n1041_ = ~new_n1040_;
  assign new_n1042_ = shift0 & a39;
  assign new_n1043_ = ~new_n1042_;
  assign new_n1044_ = new_n1043_ & new_n279_;
  assign new_n1045_ = ~new_n1044_;
  assign new_n1046_ = new_n269_ & a38;
  assign new_n1047_ = ~new_n1046_;
  assign new_n1048_ = new_n1047_ & shift1;
  assign new_n1049_ = ~new_n1048_;
  assign new_n1050_ = new_n1049_ & new_n1045_;
  assign new_n1051_ = ~new_n1050_;
  assign new_n1052_ = shift0 & a37;
  assign new_n1053_ = new_n1052_ & shift1;
  assign new_n1054_ = ~new_n1053_;
  assign new_n1055_ = new_n269_ & a40;
  assign new_n1056_ = new_n1055_ & new_n279_;
  assign new_n1057_ = ~new_n1056_;
  assign new_n1058_ = new_n1057_ & new_n1054_;
  assign new_n1059_ = new_n1058_ & new_n1051_;
  assign new_n1060_ = ~new_n1059_;
  assign new_n1061_ = new_n1060_ & new_n342_;
  assign new_n1062_ = ~new_n1061_;
  assign new_n1063_ = new_n1062_ & new_n1041_;
  assign new_n1064_ = new_n1063_ & new_n1018_;
  assign new_n1065_ = ~new_n1064_;
  assign new_n1066_ = new_n1065_ & new_n669_;
  assign new_n1067_ = ~new_n1066_;
  assign new_n1068_ = new_n1067_ & new_n971_;
  assign new_n1069_ = new_n1068_ & new_n873_;
  assign new_n1070_ = ~new_n1069_;
  assign new_n1071_ = new_n1070_ & shift6;
  assign new_n1072_ = ~new_n1071_;
  assign new_n1073_ = new_n1072_ & new_n676_;
  assign ores0 = ~new_n1073_;
  assign new_n1075_ = shift0 & a80;
  assign new_n1076_ = ~new_n1075_;
  assign new_n1077_ = new_n1076_ & new_n279_;
  assign new_n1078_ = ~new_n1077_;
  assign new_n1079_ = new_n269_ & a79;
  assign new_n1080_ = ~new_n1079_;
  assign new_n1081_ = new_n1080_ & shift1;
  assign new_n1082_ = ~new_n1081_;
  assign new_n1083_ = new_n1082_ & new_n1078_;
  assign new_n1084_ = ~new_n1083_;
  assign new_n1085_ = shift0 & a78;
  assign new_n1086_ = new_n1085_ & shift1;
  assign new_n1087_ = ~new_n1086_;
  assign new_n1088_ = new_n269_ & a81;
  assign new_n1089_ = new_n1088_ & new_n279_;
  assign new_n1090_ = ~new_n1089_;
  assign new_n1091_ = new_n1090_ & new_n1087_;
  assign new_n1092_ = new_n1091_ & new_n1084_;
  assign new_n1093_ = ~new_n1092_;
  assign new_n1094_ = new_n1093_ & new_n267_;
  assign new_n1095_ = ~new_n1094_;
  assign new_n1096_ = shift0 & a76;
  assign new_n1097_ = ~new_n1096_;
  assign new_n1098_ = new_n1097_ & new_n279_;
  assign new_n1099_ = ~new_n1098_;
  assign new_n1100_ = new_n269_ & a75;
  assign new_n1101_ = ~new_n1100_;
  assign new_n1102_ = new_n1101_ & shift1;
  assign new_n1103_ = ~new_n1102_;
  assign new_n1104_ = new_n1103_ & new_n1099_;
  assign new_n1105_ = ~new_n1104_;
  assign new_n1106_ = shift0 & a74;
  assign new_n1107_ = new_n1106_ & shift1;
  assign new_n1108_ = ~new_n1107_;
  assign new_n1109_ = new_n269_ & a77;
  assign new_n1110_ = new_n1109_ & new_n279_;
  assign new_n1111_ = ~new_n1110_;
  assign new_n1112_ = new_n1111_ & new_n1108_;
  assign new_n1113_ = new_n1112_ & new_n1105_;
  assign new_n1114_ = ~new_n1113_;
  assign new_n1115_ = new_n1114_ & new_n293_;
  assign new_n1116_ = ~new_n1115_;
  assign new_n1117_ = new_n1116_ & new_n1095_;
  assign new_n1118_ = shift0 & a68;
  assign new_n1119_ = ~new_n1118_;
  assign new_n1120_ = new_n1119_ & new_n279_;
  assign new_n1121_ = ~new_n1120_;
  assign new_n1122_ = new_n269_ & a67;
  assign new_n1123_ = ~new_n1122_;
  assign new_n1124_ = new_n1123_ & shift1;
  assign new_n1125_ = ~new_n1124_;
  assign new_n1126_ = new_n1125_ & new_n1121_;
  assign new_n1127_ = ~new_n1126_;
  assign new_n1128_ = shift0 & a66;
  assign new_n1129_ = new_n1128_ & shift1;
  assign new_n1130_ = ~new_n1129_;
  assign new_n1131_ = new_n269_ & a69;
  assign new_n1132_ = new_n1131_ & new_n279_;
  assign new_n1133_ = ~new_n1132_;
  assign new_n1134_ = new_n1133_ & new_n1130_;
  assign new_n1135_ = new_n1134_ & new_n1127_;
  assign new_n1136_ = ~new_n1135_;
  assign new_n1137_ = new_n1136_ & new_n318_;
  assign new_n1138_ = ~new_n1137_;
  assign new_n1139_ = shift0 & a72;
  assign new_n1140_ = ~new_n1139_;
  assign new_n1141_ = new_n1140_ & new_n279_;
  assign new_n1142_ = ~new_n1141_;
  assign new_n1143_ = new_n269_ & a71;
  assign new_n1144_ = ~new_n1143_;
  assign new_n1145_ = new_n1144_ & shift1;
  assign new_n1146_ = ~new_n1145_;
  assign new_n1147_ = new_n1146_ & new_n1142_;
  assign new_n1148_ = ~new_n1147_;
  assign new_n1149_ = shift0 & a70;
  assign new_n1150_ = new_n1149_ & shift1;
  assign new_n1151_ = ~new_n1150_;
  assign new_n1152_ = new_n269_ & a73;
  assign new_n1153_ = new_n1152_ & new_n279_;
  assign new_n1154_ = ~new_n1153_;
  assign new_n1155_ = new_n1154_ & new_n1151_;
  assign new_n1156_ = new_n1155_ & new_n1148_;
  assign new_n1157_ = ~new_n1156_;
  assign new_n1158_ = new_n1157_ & new_n342_;
  assign new_n1159_ = ~new_n1158_;
  assign new_n1160_ = new_n1159_ & new_n1138_;
  assign new_n1161_ = new_n1160_ & new_n1117_;
  assign new_n1162_ = ~new_n1161_;
  assign new_n1163_ = new_n1162_ & new_n369_;
  assign new_n1164_ = ~new_n1163_;
  assign new_n1165_ = shift0 & a96;
  assign new_n1166_ = ~new_n1165_;
  assign new_n1167_ = new_n1166_ & new_n279_;
  assign new_n1168_ = ~new_n1167_;
  assign new_n1169_ = new_n269_ & a95;
  assign new_n1170_ = ~new_n1169_;
  assign new_n1171_ = new_n1170_ & shift1;
  assign new_n1172_ = ~new_n1171_;
  assign new_n1173_ = new_n1172_ & new_n1168_;
  assign new_n1174_ = ~new_n1173_;
  assign new_n1175_ = shift0 & a94;
  assign new_n1176_ = new_n1175_ & shift1;
  assign new_n1177_ = ~new_n1176_;
  assign new_n1178_ = new_n269_ & a97;
  assign new_n1179_ = new_n1178_ & new_n279_;
  assign new_n1180_ = ~new_n1179_;
  assign new_n1181_ = new_n1180_ & new_n1177_;
  assign new_n1182_ = new_n1181_ & new_n1174_;
  assign new_n1183_ = ~new_n1182_;
  assign new_n1184_ = new_n1183_ & new_n267_;
  assign new_n1185_ = ~new_n1184_;
  assign new_n1186_ = shift0 & a92;
  assign new_n1187_ = ~new_n1186_;
  assign new_n1188_ = new_n1187_ & new_n279_;
  assign new_n1189_ = ~new_n1188_;
  assign new_n1190_ = new_n269_ & a91;
  assign new_n1191_ = ~new_n1190_;
  assign new_n1192_ = new_n1191_ & shift1;
  assign new_n1193_ = ~new_n1192_;
  assign new_n1194_ = new_n1193_ & new_n1189_;
  assign new_n1195_ = ~new_n1194_;
  assign new_n1196_ = shift0 & a90;
  assign new_n1197_ = new_n1196_ & shift1;
  assign new_n1198_ = ~new_n1197_;
  assign new_n1199_ = new_n269_ & a93;
  assign new_n1200_ = new_n1199_ & new_n279_;
  assign new_n1201_ = ~new_n1200_;
  assign new_n1202_ = new_n1201_ & new_n1198_;
  assign new_n1203_ = new_n1202_ & new_n1195_;
  assign new_n1204_ = ~new_n1203_;
  assign new_n1205_ = new_n1204_ & new_n293_;
  assign new_n1206_ = ~new_n1205_;
  assign new_n1207_ = new_n1206_ & new_n1185_;
  assign new_n1208_ = shift0 & a84;
  assign new_n1209_ = ~new_n1208_;
  assign new_n1210_ = new_n1209_ & new_n279_;
  assign new_n1211_ = ~new_n1210_;
  assign new_n1212_ = new_n269_ & a83;
  assign new_n1213_ = ~new_n1212_;
  assign new_n1214_ = new_n1213_ & shift1;
  assign new_n1215_ = ~new_n1214_;
  assign new_n1216_ = new_n1215_ & new_n1211_;
  assign new_n1217_ = ~new_n1216_;
  assign new_n1218_ = shift0 & a82;
  assign new_n1219_ = new_n1218_ & shift1;
  assign new_n1220_ = ~new_n1219_;
  assign new_n1221_ = new_n269_ & a85;
  assign new_n1222_ = new_n1221_ & new_n279_;
  assign new_n1223_ = ~new_n1222_;
  assign new_n1224_ = new_n1223_ & new_n1220_;
  assign new_n1225_ = new_n1224_ & new_n1217_;
  assign new_n1226_ = ~new_n1225_;
  assign new_n1227_ = new_n1226_ & new_n318_;
  assign new_n1228_ = ~new_n1227_;
  assign new_n1229_ = shift0 & a88;
  assign new_n1230_ = ~new_n1229_;
  assign new_n1231_ = new_n1230_ & new_n279_;
  assign new_n1232_ = ~new_n1231_;
  assign new_n1233_ = new_n269_ & a87;
  assign new_n1234_ = ~new_n1233_;
  assign new_n1235_ = new_n1234_ & shift1;
  assign new_n1236_ = ~new_n1235_;
  assign new_n1237_ = new_n1236_ & new_n1232_;
  assign new_n1238_ = ~new_n1237_;
  assign new_n1239_ = shift0 & a86;
  assign new_n1240_ = new_n1239_ & shift1;
  assign new_n1241_ = ~new_n1240_;
  assign new_n1242_ = new_n269_ & a89;
  assign new_n1243_ = new_n1242_ & new_n279_;
  assign new_n1244_ = ~new_n1243_;
  assign new_n1245_ = new_n1244_ & new_n1241_;
  assign new_n1246_ = new_n1245_ & new_n1238_;
  assign new_n1247_ = ~new_n1246_;
  assign new_n1248_ = new_n1247_ & new_n342_;
  assign new_n1249_ = ~new_n1248_;
  assign new_n1250_ = new_n1249_ & new_n1228_;
  assign new_n1251_ = new_n1250_ & new_n1207_;
  assign new_n1252_ = ~new_n1251_;
  assign new_n1253_ = new_n1252_ & new_n469_;
  assign new_n1254_ = ~new_n1253_;
  assign new_n1255_ = new_n1254_ & new_n1164_;
  assign new_n1256_ = shift0 & a0;
  assign new_n1257_ = ~new_n1256_;
  assign new_n1258_ = new_n1257_ & new_n279_;
  assign new_n1259_ = ~new_n1258_;
  assign new_n1260_ = new_n269_ & a127;
  assign new_n1261_ = ~new_n1260_;
  assign new_n1262_ = new_n1261_ & shift1;
  assign new_n1263_ = ~new_n1262_;
  assign new_n1264_ = new_n1263_ & new_n1259_;
  assign new_n1265_ = ~new_n1264_;
  assign new_n1266_ = shift0 & a126;
  assign new_n1267_ = new_n1266_ & shift1;
  assign new_n1268_ = ~new_n1267_;
  assign new_n1269_ = new_n269_ & a1;
  assign new_n1270_ = new_n1269_ & new_n279_;
  assign new_n1271_ = ~new_n1270_;
  assign new_n1272_ = new_n1271_ & new_n1268_;
  assign new_n1273_ = new_n1272_ & new_n1265_;
  assign new_n1274_ = ~new_n1273_;
  assign new_n1275_ = new_n1274_ & new_n267_;
  assign new_n1276_ = ~new_n1275_;
  assign new_n1277_ = shift0 & a124;
  assign new_n1278_ = ~new_n1277_;
  assign new_n1279_ = new_n1278_ & new_n279_;
  assign new_n1280_ = ~new_n1279_;
  assign new_n1281_ = new_n269_ & a123;
  assign new_n1282_ = ~new_n1281_;
  assign new_n1283_ = new_n1282_ & shift1;
  assign new_n1284_ = ~new_n1283_;
  assign new_n1285_ = new_n1284_ & new_n1280_;
  assign new_n1286_ = ~new_n1285_;
  assign new_n1287_ = shift0 & a122;
  assign new_n1288_ = new_n1287_ & shift1;
  assign new_n1289_ = ~new_n1288_;
  assign new_n1290_ = new_n269_ & a125;
  assign new_n1291_ = new_n1290_ & new_n279_;
  assign new_n1292_ = ~new_n1291_;
  assign new_n1293_ = new_n1292_ & new_n1289_;
  assign new_n1294_ = new_n1293_ & new_n1286_;
  assign new_n1295_ = ~new_n1294_;
  assign new_n1296_ = new_n1295_ & new_n293_;
  assign new_n1297_ = ~new_n1296_;
  assign new_n1298_ = new_n1297_ & new_n1276_;
  assign new_n1299_ = shift0 & a116;
  assign new_n1300_ = ~new_n1299_;
  assign new_n1301_ = new_n1300_ & new_n279_;
  assign new_n1302_ = ~new_n1301_;
  assign new_n1303_ = new_n269_ & a115;
  assign new_n1304_ = ~new_n1303_;
  assign new_n1305_ = new_n1304_ & shift1;
  assign new_n1306_ = ~new_n1305_;
  assign new_n1307_ = new_n1306_ & new_n1302_;
  assign new_n1308_ = ~new_n1307_;
  assign new_n1309_ = shift0 & a114;
  assign new_n1310_ = new_n1309_ & shift1;
  assign new_n1311_ = ~new_n1310_;
  assign new_n1312_ = new_n269_ & a117;
  assign new_n1313_ = new_n1312_ & new_n279_;
  assign new_n1314_ = ~new_n1313_;
  assign new_n1315_ = new_n1314_ & new_n1311_;
  assign new_n1316_ = new_n1315_ & new_n1308_;
  assign new_n1317_ = ~new_n1316_;
  assign new_n1318_ = new_n1317_ & new_n318_;
  assign new_n1319_ = ~new_n1318_;
  assign new_n1320_ = shift0 & a120;
  assign new_n1321_ = ~new_n1320_;
  assign new_n1322_ = new_n1321_ & new_n279_;
  assign new_n1323_ = ~new_n1322_;
  assign new_n1324_ = new_n269_ & a119;
  assign new_n1325_ = ~new_n1324_;
  assign new_n1326_ = new_n1325_ & shift1;
  assign new_n1327_ = ~new_n1326_;
  assign new_n1328_ = new_n1327_ & new_n1323_;
  assign new_n1329_ = ~new_n1328_;
  assign new_n1330_ = shift0 & a118;
  assign new_n1331_ = new_n1330_ & shift1;
  assign new_n1332_ = ~new_n1331_;
  assign new_n1333_ = new_n269_ & a121;
  assign new_n1334_ = new_n1333_ & new_n279_;
  assign new_n1335_ = ~new_n1334_;
  assign new_n1336_ = new_n1335_ & new_n1332_;
  assign new_n1337_ = new_n1336_ & new_n1329_;
  assign new_n1338_ = ~new_n1337_;
  assign new_n1339_ = new_n1338_ & new_n342_;
  assign new_n1340_ = ~new_n1339_;
  assign new_n1341_ = new_n1340_ & new_n1319_;
  assign new_n1342_ = new_n1341_ & new_n1298_;
  assign new_n1343_ = ~new_n1342_;
  assign new_n1344_ = new_n1343_ & new_n570_;
  assign new_n1345_ = ~new_n1344_;
  assign new_n1346_ = shift0 & a112;
  assign new_n1347_ = ~new_n1346_;
  assign new_n1348_ = new_n1347_ & new_n279_;
  assign new_n1349_ = ~new_n1348_;
  assign new_n1350_ = new_n269_ & a111;
  assign new_n1351_ = ~new_n1350_;
  assign new_n1352_ = new_n1351_ & shift1;
  assign new_n1353_ = ~new_n1352_;
  assign new_n1354_ = new_n1353_ & new_n1349_;
  assign new_n1355_ = ~new_n1354_;
  assign new_n1356_ = shift0 & a110;
  assign new_n1357_ = new_n1356_ & shift1;
  assign new_n1358_ = ~new_n1357_;
  assign new_n1359_ = new_n269_ & a113;
  assign new_n1360_ = new_n1359_ & new_n279_;
  assign new_n1361_ = ~new_n1360_;
  assign new_n1362_ = new_n1361_ & new_n1358_;
  assign new_n1363_ = new_n1362_ & new_n1355_;
  assign new_n1364_ = ~new_n1363_;
  assign new_n1365_ = new_n1364_ & new_n267_;
  assign new_n1366_ = ~new_n1365_;
  assign new_n1367_ = shift0 & a108;
  assign new_n1368_ = ~new_n1367_;
  assign new_n1369_ = new_n1368_ & new_n279_;
  assign new_n1370_ = ~new_n1369_;
  assign new_n1371_ = new_n269_ & a107;
  assign new_n1372_ = ~new_n1371_;
  assign new_n1373_ = new_n1372_ & shift1;
  assign new_n1374_ = ~new_n1373_;
  assign new_n1375_ = new_n1374_ & new_n1370_;
  assign new_n1376_ = ~new_n1375_;
  assign new_n1377_ = shift0 & a106;
  assign new_n1378_ = new_n1377_ & shift1;
  assign new_n1379_ = ~new_n1378_;
  assign new_n1380_ = new_n269_ & a109;
  assign new_n1381_ = new_n1380_ & new_n279_;
  assign new_n1382_ = ~new_n1381_;
  assign new_n1383_ = new_n1382_ & new_n1379_;
  assign new_n1384_ = new_n1383_ & new_n1376_;
  assign new_n1385_ = ~new_n1384_;
  assign new_n1386_ = new_n1385_ & new_n293_;
  assign new_n1387_ = ~new_n1386_;
  assign new_n1388_ = new_n1387_ & new_n1366_;
  assign new_n1389_ = shift0 & a100;
  assign new_n1390_ = ~new_n1389_;
  assign new_n1391_ = new_n1390_ & new_n279_;
  assign new_n1392_ = ~new_n1391_;
  assign new_n1393_ = new_n269_ & a99;
  assign new_n1394_ = ~new_n1393_;
  assign new_n1395_ = new_n1394_ & shift1;
  assign new_n1396_ = ~new_n1395_;
  assign new_n1397_ = new_n1396_ & new_n1392_;
  assign new_n1398_ = ~new_n1397_;
  assign new_n1399_ = shift0 & a98;
  assign new_n1400_ = new_n1399_ & shift1;
  assign new_n1401_ = ~new_n1400_;
  assign new_n1402_ = new_n269_ & a101;
  assign new_n1403_ = new_n1402_ & new_n279_;
  assign new_n1404_ = ~new_n1403_;
  assign new_n1405_ = new_n1404_ & new_n1401_;
  assign new_n1406_ = new_n1405_ & new_n1398_;
  assign new_n1407_ = ~new_n1406_;
  assign new_n1408_ = new_n1407_ & new_n318_;
  assign new_n1409_ = ~new_n1408_;
  assign new_n1410_ = shift0 & a104;
  assign new_n1411_ = ~new_n1410_;
  assign new_n1412_ = new_n1411_ & new_n279_;
  assign new_n1413_ = ~new_n1412_;
  assign new_n1414_ = new_n269_ & a103;
  assign new_n1415_ = ~new_n1414_;
  assign new_n1416_ = new_n1415_ & shift1;
  assign new_n1417_ = ~new_n1416_;
  assign new_n1418_ = new_n1417_ & new_n1413_;
  assign new_n1419_ = ~new_n1418_;
  assign new_n1420_ = shift0 & a102;
  assign new_n1421_ = new_n1420_ & shift1;
  assign new_n1422_ = ~new_n1421_;
  assign new_n1423_ = new_n269_ & a105;
  assign new_n1424_ = new_n1423_ & new_n279_;
  assign new_n1425_ = ~new_n1424_;
  assign new_n1426_ = new_n1425_ & new_n1422_;
  assign new_n1427_ = new_n1426_ & new_n1419_;
  assign new_n1428_ = ~new_n1427_;
  assign new_n1429_ = new_n1428_ & new_n342_;
  assign new_n1430_ = ~new_n1429_;
  assign new_n1431_ = new_n1430_ & new_n1409_;
  assign new_n1432_ = new_n1431_ & new_n1388_;
  assign new_n1433_ = ~new_n1432_;
  assign new_n1434_ = new_n1433_ & new_n669_;
  assign new_n1435_ = ~new_n1434_;
  assign new_n1436_ = new_n1435_ & new_n1345_;
  assign new_n1437_ = new_n1436_ & new_n1255_;
  assign new_n1438_ = ~new_n1437_;
  assign new_n1439_ = new_n1438_ & new_n264_;
  assign new_n1440_ = ~new_n1439_;
  assign new_n1441_ = shift0 & a64;
  assign new_n1442_ = ~new_n1441_;
  assign new_n1443_ = new_n1442_ & new_n279_;
  assign new_n1444_ = ~new_n1443_;
  assign new_n1445_ = new_n269_ & a63;
  assign new_n1446_ = ~new_n1445_;
  assign new_n1447_ = new_n1446_ & shift1;
  assign new_n1448_ = ~new_n1447_;
  assign new_n1449_ = new_n1448_ & new_n1444_;
  assign new_n1450_ = ~new_n1449_;
  assign new_n1451_ = shift0 & a62;
  assign new_n1452_ = new_n1451_ & shift1;
  assign new_n1453_ = ~new_n1452_;
  assign new_n1454_ = new_n269_ & a65;
  assign new_n1455_ = new_n1454_ & new_n279_;
  assign new_n1456_ = ~new_n1455_;
  assign new_n1457_ = new_n1456_ & new_n1453_;
  assign new_n1458_ = new_n1457_ & new_n1450_;
  assign new_n1459_ = ~new_n1458_;
  assign new_n1460_ = new_n1459_ & new_n267_;
  assign new_n1461_ = ~new_n1460_;
  assign new_n1462_ = shift0 & a60;
  assign new_n1463_ = ~new_n1462_;
  assign new_n1464_ = new_n1463_ & new_n279_;
  assign new_n1465_ = ~new_n1464_;
  assign new_n1466_ = new_n269_ & a59;
  assign new_n1467_ = ~new_n1466_;
  assign new_n1468_ = new_n1467_ & shift1;
  assign new_n1469_ = ~new_n1468_;
  assign new_n1470_ = new_n1469_ & new_n1465_;
  assign new_n1471_ = ~new_n1470_;
  assign new_n1472_ = shift0 & a58;
  assign new_n1473_ = new_n1472_ & shift1;
  assign new_n1474_ = ~new_n1473_;
  assign new_n1475_ = new_n269_ & a61;
  assign new_n1476_ = new_n1475_ & new_n279_;
  assign new_n1477_ = ~new_n1476_;
  assign new_n1478_ = new_n1477_ & new_n1474_;
  assign new_n1479_ = new_n1478_ & new_n1471_;
  assign new_n1480_ = ~new_n1479_;
  assign new_n1481_ = new_n1480_ & new_n293_;
  assign new_n1482_ = ~new_n1481_;
  assign new_n1483_ = new_n1482_ & new_n1461_;
  assign new_n1484_ = shift0 & a52;
  assign new_n1485_ = ~new_n1484_;
  assign new_n1486_ = new_n1485_ & new_n279_;
  assign new_n1487_ = ~new_n1486_;
  assign new_n1488_ = new_n269_ & a51;
  assign new_n1489_ = ~new_n1488_;
  assign new_n1490_ = new_n1489_ & shift1;
  assign new_n1491_ = ~new_n1490_;
  assign new_n1492_ = new_n1491_ & new_n1487_;
  assign new_n1493_ = ~new_n1492_;
  assign new_n1494_ = shift0 & a50;
  assign new_n1495_ = new_n1494_ & shift1;
  assign new_n1496_ = ~new_n1495_;
  assign new_n1497_ = new_n269_ & a53;
  assign new_n1498_ = new_n1497_ & new_n279_;
  assign new_n1499_ = ~new_n1498_;
  assign new_n1500_ = new_n1499_ & new_n1496_;
  assign new_n1501_ = new_n1500_ & new_n1493_;
  assign new_n1502_ = ~new_n1501_;
  assign new_n1503_ = new_n1502_ & new_n318_;
  assign new_n1504_ = ~new_n1503_;
  assign new_n1505_ = shift0 & a56;
  assign new_n1506_ = ~new_n1505_;
  assign new_n1507_ = new_n1506_ & new_n279_;
  assign new_n1508_ = ~new_n1507_;
  assign new_n1509_ = new_n269_ & a55;
  assign new_n1510_ = ~new_n1509_;
  assign new_n1511_ = new_n1510_ & shift1;
  assign new_n1512_ = ~new_n1511_;
  assign new_n1513_ = new_n1512_ & new_n1508_;
  assign new_n1514_ = ~new_n1513_;
  assign new_n1515_ = shift0 & a54;
  assign new_n1516_ = new_n1515_ & shift1;
  assign new_n1517_ = ~new_n1516_;
  assign new_n1518_ = new_n269_ & a57;
  assign new_n1519_ = new_n1518_ & new_n279_;
  assign new_n1520_ = ~new_n1519_;
  assign new_n1521_ = new_n1520_ & new_n1517_;
  assign new_n1522_ = new_n1521_ & new_n1514_;
  assign new_n1523_ = ~new_n1522_;
  assign new_n1524_ = new_n1523_ & new_n342_;
  assign new_n1525_ = ~new_n1524_;
  assign new_n1526_ = new_n1525_ & new_n1504_;
  assign new_n1527_ = new_n1526_ & new_n1483_;
  assign new_n1528_ = ~new_n1527_;
  assign new_n1529_ = new_n1528_ & new_n570_;
  assign new_n1530_ = ~new_n1529_;
  assign new_n1531_ = shift0 & a16;
  assign new_n1532_ = ~new_n1531_;
  assign new_n1533_ = new_n1532_ & new_n279_;
  assign new_n1534_ = ~new_n1533_;
  assign new_n1535_ = new_n269_ & a15;
  assign new_n1536_ = ~new_n1535_;
  assign new_n1537_ = new_n1536_ & shift1;
  assign new_n1538_ = ~new_n1537_;
  assign new_n1539_ = new_n1538_ & new_n1534_;
  assign new_n1540_ = ~new_n1539_;
  assign new_n1541_ = shift0 & a14;
  assign new_n1542_ = new_n1541_ & shift1;
  assign new_n1543_ = ~new_n1542_;
  assign new_n1544_ = new_n269_ & a17;
  assign new_n1545_ = new_n1544_ & new_n279_;
  assign new_n1546_ = ~new_n1545_;
  assign new_n1547_ = new_n1546_ & new_n1543_;
  assign new_n1548_ = new_n1547_ & new_n1540_;
  assign new_n1549_ = ~new_n1548_;
  assign new_n1550_ = new_n1549_ & new_n267_;
  assign new_n1551_ = ~new_n1550_;
  assign new_n1552_ = shift0 & a12;
  assign new_n1553_ = ~new_n1552_;
  assign new_n1554_ = new_n1553_ & new_n279_;
  assign new_n1555_ = ~new_n1554_;
  assign new_n1556_ = new_n269_ & a11;
  assign new_n1557_ = ~new_n1556_;
  assign new_n1558_ = new_n1557_ & shift1;
  assign new_n1559_ = ~new_n1558_;
  assign new_n1560_ = new_n1559_ & new_n1555_;
  assign new_n1561_ = ~new_n1560_;
  assign new_n1562_ = shift0 & a10;
  assign new_n1563_ = new_n1562_ & shift1;
  assign new_n1564_ = ~new_n1563_;
  assign new_n1565_ = new_n269_ & a13;
  assign new_n1566_ = new_n1565_ & new_n279_;
  assign new_n1567_ = ~new_n1566_;
  assign new_n1568_ = new_n1567_ & new_n1564_;
  assign new_n1569_ = new_n1568_ & new_n1561_;
  assign new_n1570_ = ~new_n1569_;
  assign new_n1571_ = new_n1570_ & new_n293_;
  assign new_n1572_ = ~new_n1571_;
  assign new_n1573_ = new_n1572_ & new_n1551_;
  assign new_n1574_ = shift0 & a4;
  assign new_n1575_ = ~new_n1574_;
  assign new_n1576_ = new_n1575_ & new_n279_;
  assign new_n1577_ = ~new_n1576_;
  assign new_n1578_ = new_n269_ & a3;
  assign new_n1579_ = ~new_n1578_;
  assign new_n1580_ = new_n1579_ & shift1;
  assign new_n1581_ = ~new_n1580_;
  assign new_n1582_ = new_n1581_ & new_n1577_;
  assign new_n1583_ = ~new_n1582_;
  assign new_n1584_ = shift0 & a2;
  assign new_n1585_ = new_n1584_ & shift1;
  assign new_n1586_ = ~new_n1585_;
  assign new_n1587_ = new_n269_ & a5;
  assign new_n1588_ = new_n1587_ & new_n279_;
  assign new_n1589_ = ~new_n1588_;
  assign new_n1590_ = new_n1589_ & new_n1586_;
  assign new_n1591_ = new_n1590_ & new_n1583_;
  assign new_n1592_ = ~new_n1591_;
  assign new_n1593_ = new_n1592_ & new_n318_;
  assign new_n1594_ = ~new_n1593_;
  assign new_n1595_ = shift0 & a8;
  assign new_n1596_ = ~new_n1595_;
  assign new_n1597_ = new_n1596_ & new_n279_;
  assign new_n1598_ = ~new_n1597_;
  assign new_n1599_ = new_n269_ & a7;
  assign new_n1600_ = ~new_n1599_;
  assign new_n1601_ = new_n1600_ & shift1;
  assign new_n1602_ = ~new_n1601_;
  assign new_n1603_ = new_n1602_ & new_n1598_;
  assign new_n1604_ = ~new_n1603_;
  assign new_n1605_ = shift0 & a6;
  assign new_n1606_ = new_n1605_ & shift1;
  assign new_n1607_ = ~new_n1606_;
  assign new_n1608_ = new_n269_ & a9;
  assign new_n1609_ = new_n1608_ & new_n279_;
  assign new_n1610_ = ~new_n1609_;
  assign new_n1611_ = new_n1610_ & new_n1607_;
  assign new_n1612_ = new_n1611_ & new_n1604_;
  assign new_n1613_ = ~new_n1612_;
  assign new_n1614_ = new_n1613_ & new_n342_;
  assign new_n1615_ = ~new_n1614_;
  assign new_n1616_ = new_n1615_ & new_n1594_;
  assign new_n1617_ = new_n1616_ & new_n1573_;
  assign new_n1618_ = ~new_n1617_;
  assign new_n1619_ = new_n1618_ & new_n369_;
  assign new_n1620_ = ~new_n1619_;
  assign new_n1621_ = new_n1620_ & new_n1530_;
  assign new_n1622_ = shift0 & a48;
  assign new_n1623_ = ~new_n1622_;
  assign new_n1624_ = new_n1623_ & new_n279_;
  assign new_n1625_ = ~new_n1624_;
  assign new_n1626_ = new_n269_ & a47;
  assign new_n1627_ = ~new_n1626_;
  assign new_n1628_ = new_n1627_ & shift1;
  assign new_n1629_ = ~new_n1628_;
  assign new_n1630_ = new_n1629_ & new_n1625_;
  assign new_n1631_ = ~new_n1630_;
  assign new_n1632_ = shift0 & a46;
  assign new_n1633_ = new_n1632_ & shift1;
  assign new_n1634_ = ~new_n1633_;
  assign new_n1635_ = new_n269_ & a49;
  assign new_n1636_ = new_n1635_ & new_n279_;
  assign new_n1637_ = ~new_n1636_;
  assign new_n1638_ = new_n1637_ & new_n1634_;
  assign new_n1639_ = new_n1638_ & new_n1631_;
  assign new_n1640_ = ~new_n1639_;
  assign new_n1641_ = new_n1640_ & new_n267_;
  assign new_n1642_ = ~new_n1641_;
  assign new_n1643_ = shift0 & a42;
  assign new_n1644_ = ~new_n1643_;
  assign new_n1645_ = new_n269_ & a43;
  assign new_n1646_ = ~new_n1645_;
  assign new_n1647_ = new_n1646_ & new_n1644_;
  assign new_n1648_ = ~new_n1647_;
  assign new_n1649_ = new_n1648_ & shift1;
  assign new_n1650_ = ~new_n1649_;
  assign new_n1651_ = shift0 & new_n1008_;
  assign new_n1652_ = ~new_n1651_;
  assign new_n1653_ = new_n269_ & new_n975_;
  assign new_n1654_ = ~new_n1653_;
  assign new_n1655_ = new_n1654_ & new_n1652_;
  assign new_n1656_ = new_n1655_ & new_n279_;
  assign new_n1657_ = ~new_n1656_;
  assign new_n1658_ = new_n1657_ & new_n1650_;
  assign new_n1659_ = ~new_n1658_;
  assign new_n1660_ = new_n1659_ & new_n293_;
  assign new_n1661_ = ~new_n1660_;
  assign new_n1662_ = new_n1661_ & new_n1642_;
  assign new_n1663_ = shift0 & a36;
  assign new_n1664_ = ~new_n1663_;
  assign new_n1665_ = new_n1664_ & new_n279_;
  assign new_n1666_ = ~new_n1665_;
  assign new_n1667_ = new_n269_ & a35;
  assign new_n1668_ = ~new_n1667_;
  assign new_n1669_ = new_n1668_ & shift1;
  assign new_n1670_ = ~new_n1669_;
  assign new_n1671_ = new_n1670_ & new_n1666_;
  assign new_n1672_ = ~new_n1671_;
  assign new_n1673_ = shift0 & a34;
  assign new_n1674_ = new_n1673_ & shift1;
  assign new_n1675_ = ~new_n1674_;
  assign new_n1676_ = new_n269_ & a37;
  assign new_n1677_ = new_n1676_ & new_n279_;
  assign new_n1678_ = ~new_n1677_;
  assign new_n1679_ = new_n1678_ & new_n1675_;
  assign new_n1680_ = new_n1679_ & new_n1672_;
  assign new_n1681_ = ~new_n1680_;
  assign new_n1682_ = new_n1681_ & new_n318_;
  assign new_n1683_ = ~new_n1682_;
  assign new_n1684_ = new_n269_ & a41;
  assign new_n1685_ = ~new_n1684_;
  assign new_n1686_ = shift0 & a40;
  assign new_n1687_ = ~new_n1686_;
  assign new_n1688_ = new_n1687_ & new_n1685_;
  assign new_n1689_ = ~new_n1688_;
  assign new_n1690_ = new_n1689_ & new_n279_;
  assign new_n1691_ = ~new_n1690_;
  assign new_n1692_ = new_n269_ & a39;
  assign new_n1693_ = ~new_n1692_;
  assign new_n1694_ = shift0 & a38;
  assign new_n1695_ = ~new_n1694_;
  assign new_n1696_ = new_n1695_ & new_n1693_;
  assign new_n1697_ = ~new_n1696_;
  assign new_n1698_ = new_n1697_ & shift1;
  assign new_n1699_ = ~new_n1698_;
  assign new_n1700_ = new_n1699_ & new_n1691_;
  assign new_n1701_ = ~new_n1700_;
  assign new_n1702_ = new_n1701_ & new_n342_;
  assign new_n1703_ = ~new_n1702_;
  assign new_n1704_ = new_n1703_ & new_n1683_;
  assign new_n1705_ = new_n1704_ & new_n1662_;
  assign new_n1706_ = ~new_n1705_;
  assign new_n1707_ = new_n1706_ & new_n669_;
  assign new_n1708_ = ~new_n1707_;
  assign new_n1709_ = shift0 & a32;
  assign new_n1710_ = ~new_n1709_;
  assign new_n1711_ = new_n1710_ & new_n279_;
  assign new_n1712_ = ~new_n1711_;
  assign new_n1713_ = new_n269_ & a31;
  assign new_n1714_ = ~new_n1713_;
  assign new_n1715_ = new_n1714_ & shift1;
  assign new_n1716_ = ~new_n1715_;
  assign new_n1717_ = new_n1716_ & new_n1712_;
  assign new_n1718_ = ~new_n1717_;
  assign new_n1719_ = shift0 & a30;
  assign new_n1720_ = new_n1719_ & shift1;
  assign new_n1721_ = ~new_n1720_;
  assign new_n1722_ = new_n269_ & a33;
  assign new_n1723_ = new_n1722_ & new_n279_;
  assign new_n1724_ = ~new_n1723_;
  assign new_n1725_ = new_n1724_ & new_n1721_;
  assign new_n1726_ = new_n1725_ & new_n1718_;
  assign new_n1727_ = ~new_n1726_;
  assign new_n1728_ = new_n1727_ & new_n267_;
  assign new_n1729_ = ~new_n1728_;
  assign new_n1730_ = shift0 & a28;
  assign new_n1731_ = ~new_n1730_;
  assign new_n1732_ = new_n1731_ & new_n279_;
  assign new_n1733_ = ~new_n1732_;
  assign new_n1734_ = new_n269_ & a27;
  assign new_n1735_ = ~new_n1734_;
  assign new_n1736_ = new_n1735_ & shift1;
  assign new_n1737_ = ~new_n1736_;
  assign new_n1738_ = new_n1737_ & new_n1733_;
  assign new_n1739_ = ~new_n1738_;
  assign new_n1740_ = shift0 & a26;
  assign new_n1741_ = new_n1740_ & shift1;
  assign new_n1742_ = ~new_n1741_;
  assign new_n1743_ = new_n269_ & a29;
  assign new_n1744_ = new_n1743_ & new_n279_;
  assign new_n1745_ = ~new_n1744_;
  assign new_n1746_ = new_n1745_ & new_n1742_;
  assign new_n1747_ = new_n1746_ & new_n1739_;
  assign new_n1748_ = ~new_n1747_;
  assign new_n1749_ = new_n1748_ & new_n293_;
  assign new_n1750_ = ~new_n1749_;
  assign new_n1751_ = new_n1750_ & new_n1729_;
  assign new_n1752_ = shift0 & a20;
  assign new_n1753_ = ~new_n1752_;
  assign new_n1754_ = new_n1753_ & new_n279_;
  assign new_n1755_ = ~new_n1754_;
  assign new_n1756_ = new_n269_ & a19;
  assign new_n1757_ = ~new_n1756_;
  assign new_n1758_ = new_n1757_ & shift1;
  assign new_n1759_ = ~new_n1758_;
  assign new_n1760_ = new_n1759_ & new_n1755_;
  assign new_n1761_ = ~new_n1760_;
  assign new_n1762_ = shift0 & a18;
  assign new_n1763_ = new_n1762_ & shift1;
  assign new_n1764_ = ~new_n1763_;
  assign new_n1765_ = new_n269_ & a21;
  assign new_n1766_ = new_n1765_ & new_n279_;
  assign new_n1767_ = ~new_n1766_;
  assign new_n1768_ = new_n1767_ & new_n1764_;
  assign new_n1769_ = new_n1768_ & new_n1761_;
  assign new_n1770_ = ~new_n1769_;
  assign new_n1771_ = new_n1770_ & new_n318_;
  assign new_n1772_ = ~new_n1771_;
  assign new_n1773_ = shift0 & a24;
  assign new_n1774_ = ~new_n1773_;
  assign new_n1775_ = new_n1774_ & new_n279_;
  assign new_n1776_ = ~new_n1775_;
  assign new_n1777_ = new_n269_ & a23;
  assign new_n1778_ = ~new_n1777_;
  assign new_n1779_ = new_n1778_ & shift1;
  assign new_n1780_ = ~new_n1779_;
  assign new_n1781_ = new_n1780_ & new_n1776_;
  assign new_n1782_ = ~new_n1781_;
  assign new_n1783_ = shift0 & a22;
  assign new_n1784_ = new_n1783_ & shift1;
  assign new_n1785_ = ~new_n1784_;
  assign new_n1786_ = new_n269_ & a25;
  assign new_n1787_ = new_n1786_ & new_n279_;
  assign new_n1788_ = ~new_n1787_;
  assign new_n1789_ = new_n1788_ & new_n1785_;
  assign new_n1790_ = new_n1789_ & new_n1782_;
  assign new_n1791_ = ~new_n1790_;
  assign new_n1792_ = new_n1791_ & new_n342_;
  assign new_n1793_ = ~new_n1792_;
  assign new_n1794_ = new_n1793_ & new_n1772_;
  assign new_n1795_ = new_n1794_ & new_n1751_;
  assign new_n1796_ = ~new_n1795_;
  assign new_n1797_ = new_n1796_ & new_n469_;
  assign new_n1798_ = ~new_n1797_;
  assign new_n1799_ = new_n1798_ & new_n1708_;
  assign new_n1800_ = new_n1799_ & new_n1621_;
  assign new_n1801_ = ~new_n1800_;
  assign new_n1802_ = new_n1801_ & shift6;
  assign new_n1803_ = ~new_n1802_;
  assign new_n1804_ = new_n1803_ & new_n1440_;
  assign ores1 = ~new_n1804_;
  assign new_n1806_ = new_n287_ & shift1;
  assign new_n1807_ = ~new_n1806_;
  assign new_n1808_ = new_n426_ & new_n279_;
  assign new_n1809_ = ~new_n1808_;
  assign new_n1810_ = new_n1809_ & new_n1807_;
  assign new_n1811_ = new_n1810_ & new_n267_;
  assign new_n1812_ = ~new_n1811_;
  assign new_n1813_ = new_n311_ & shift1;
  assign new_n1814_ = ~new_n1813_;
  assign new_n1815_ = new_n276_ & new_n279_;
  assign new_n1816_ = ~new_n1815_;
  assign new_n1817_ = new_n1816_ & new_n1814_;
  assign new_n1818_ = new_n1817_ & new_n293_;
  assign new_n1819_ = ~new_n1818_;
  assign new_n1820_ = new_n1819_ & new_n1812_;
  assign new_n1821_ = new_n336_ & shift1;
  assign new_n1822_ = ~new_n1821_;
  assign new_n1823_ = new_n350_ & new_n279_;
  assign new_n1824_ = ~new_n1823_;
  assign new_n1825_ = new_n1824_ & new_n1822_;
  assign new_n1826_ = new_n1825_ & new_n318_;
  assign new_n1827_ = ~new_n1826_;
  assign new_n1828_ = new_n360_ & shift1;
  assign new_n1829_ = ~new_n1828_;
  assign new_n1830_ = new_n301_ & new_n279_;
  assign new_n1831_ = ~new_n1830_;
  assign new_n1832_ = new_n1831_ & new_n1829_;
  assign new_n1833_ = new_n1832_ & new_n342_;
  assign new_n1834_ = ~new_n1833_;
  assign new_n1835_ = new_n1834_ & new_n1827_;
  assign new_n1836_ = new_n1835_ & new_n1820_;
  assign new_n1837_ = ~new_n1836_;
  assign new_n1838_ = new_n1837_ & new_n369_;
  assign new_n1839_ = ~new_n1838_;
  assign new_n1840_ = new_n389_ & shift1;
  assign new_n1841_ = ~new_n1840_;
  assign new_n1842_ = new_n627_ & new_n279_;
  assign new_n1843_ = ~new_n1842_;
  assign new_n1844_ = new_n1843_ & new_n1841_;
  assign new_n1845_ = new_n1844_ & new_n267_;
  assign new_n1846_ = ~new_n1845_;
  assign new_n1847_ = new_n412_ & shift1;
  assign new_n1848_ = ~new_n1847_;
  assign new_n1849_ = new_n379_ & new_n279_;
  assign new_n1850_ = ~new_n1849_;
  assign new_n1851_ = new_n1850_ & new_n1848_;
  assign new_n1852_ = new_n1851_ & new_n293_;
  assign new_n1853_ = ~new_n1852_;
  assign new_n1854_ = new_n1853_ & new_n1846_;
  assign new_n1855_ = new_n436_ & shift1;
  assign new_n1856_ = ~new_n1855_;
  assign new_n1857_ = new_n449_ & new_n279_;
  assign new_n1858_ = ~new_n1857_;
  assign new_n1859_ = new_n1858_ & new_n1856_;
  assign new_n1860_ = new_n1859_ & new_n318_;
  assign new_n1861_ = ~new_n1860_;
  assign new_n1862_ = new_n459_ & shift1;
  assign new_n1863_ = ~new_n1862_;
  assign new_n1864_ = new_n402_ & new_n279_;
  assign new_n1865_ = ~new_n1864_;
  assign new_n1866_ = new_n1865_ & new_n1863_;
  assign new_n1867_ = new_n1866_ & new_n342_;
  assign new_n1868_ = ~new_n1867_;
  assign new_n1869_ = new_n1868_ & new_n1861_;
  assign new_n1870_ = new_n1869_ & new_n1854_;
  assign new_n1871_ = ~new_n1870_;
  assign new_n1872_ = new_n1871_ & new_n469_;
  assign new_n1873_ = ~new_n1872_;
  assign new_n1874_ = new_n1873_ & new_n1839_;
  assign new_n1875_ = new_n490_ & shift1;
  assign new_n1876_ = ~new_n1875_;
  assign new_n1877_ = new_n731_ & new_n279_;
  assign new_n1878_ = ~new_n1877_;
  assign new_n1879_ = new_n1878_ & new_n1876_;
  assign new_n1880_ = new_n1879_ & new_n267_;
  assign new_n1881_ = ~new_n1880_;
  assign new_n1882_ = new_n513_ & shift1;
  assign new_n1883_ = ~new_n1882_;
  assign new_n1884_ = new_n480_ & new_n279_;
  assign new_n1885_ = ~new_n1884_;
  assign new_n1886_ = new_n1885_ & new_n1883_;
  assign new_n1887_ = new_n1886_ & new_n293_;
  assign new_n1888_ = ~new_n1887_;
  assign new_n1889_ = new_n1888_ & new_n1881_;
  assign new_n1890_ = new_n537_ & shift1;
  assign new_n1891_ = ~new_n1890_;
  assign new_n1892_ = new_n550_ & new_n279_;
  assign new_n1893_ = ~new_n1892_;
  assign new_n1894_ = new_n1893_ & new_n1891_;
  assign new_n1895_ = new_n1894_ & new_n318_;
  assign new_n1896_ = ~new_n1895_;
  assign new_n1897_ = new_n560_ & shift1;
  assign new_n1898_ = ~new_n1897_;
  assign new_n1899_ = new_n503_ & new_n279_;
  assign new_n1900_ = ~new_n1899_;
  assign new_n1901_ = new_n1900_ & new_n1898_;
  assign new_n1902_ = new_n1901_ & new_n342_;
  assign new_n1903_ = ~new_n1902_;
  assign new_n1904_ = new_n1903_ & new_n1896_;
  assign new_n1905_ = new_n1904_ & new_n1889_;
  assign new_n1906_ = ~new_n1905_;
  assign new_n1907_ = new_n1906_ & new_n570_;
  assign new_n1908_ = ~new_n1907_;
  assign new_n1909_ = new_n590_ & shift1;
  assign new_n1910_ = ~new_n1909_;
  assign new_n1911_ = new_n527_ & new_n279_;
  assign new_n1912_ = ~new_n1911_;
  assign new_n1913_ = new_n1912_ & new_n1910_;
  assign new_n1914_ = new_n1913_ & new_n267_;
  assign new_n1915_ = ~new_n1914_;
  assign new_n1916_ = new_n613_ & shift1;
  assign new_n1917_ = ~new_n1916_;
  assign new_n1918_ = new_n580_ & new_n279_;
  assign new_n1919_ = ~new_n1918_;
  assign new_n1920_ = new_n1919_ & new_n1917_;
  assign new_n1921_ = new_n1920_ & new_n293_;
  assign new_n1922_ = ~new_n1921_;
  assign new_n1923_ = new_n1922_ & new_n1915_;
  assign new_n1924_ = new_n637_ & shift1;
  assign new_n1925_ = ~new_n1924_;
  assign new_n1926_ = new_n650_ & new_n279_;
  assign new_n1927_ = ~new_n1926_;
  assign new_n1928_ = new_n1927_ & new_n1925_;
  assign new_n1929_ = new_n1928_ & new_n318_;
  assign new_n1930_ = ~new_n1929_;
  assign new_n1931_ = new_n660_ & shift1;
  assign new_n1932_ = ~new_n1931_;
  assign new_n1933_ = new_n603_ & new_n279_;
  assign new_n1934_ = ~new_n1933_;
  assign new_n1935_ = new_n1934_ & new_n1932_;
  assign new_n1936_ = new_n1935_ & new_n342_;
  assign new_n1937_ = ~new_n1936_;
  assign new_n1938_ = new_n1937_ & new_n1930_;
  assign new_n1939_ = new_n1938_ & new_n1923_;
  assign new_n1940_ = ~new_n1939_;
  assign new_n1941_ = new_n1940_ & new_n669_;
  assign new_n1942_ = ~new_n1941_;
  assign new_n1943_ = new_n1942_ & new_n1908_;
  assign new_n1944_ = new_n1943_ & new_n1874_;
  assign new_n1945_ = ~new_n1944_;
  assign new_n1946_ = new_n1945_ & new_n264_;
  assign new_n1947_ = ~new_n1946_;
  assign new_n1948_ = new_n891_ & shift1;
  assign new_n1949_ = ~new_n1948_;
  assign new_n1950_ = new_n326_ & new_n279_;
  assign new_n1951_ = ~new_n1950_;
  assign new_n1952_ = new_n1951_ & new_n1949_;
  assign new_n1953_ = new_n1952_ & new_n267_;
  assign new_n1954_ = ~new_n1953_;
  assign new_n1955_ = new_n914_ & shift1;
  assign new_n1956_ = ~new_n1955_;
  assign new_n1957_ = new_n881_ & new_n279_;
  assign new_n1958_ = ~new_n1957_;
  assign new_n1959_ = new_n1958_ & new_n1956_;
  assign new_n1960_ = new_n1959_ & new_n293_;
  assign new_n1961_ = ~new_n1960_;
  assign new_n1962_ = new_n1961_ & new_n1954_;
  assign new_n1963_ = new_n938_ & shift1;
  assign new_n1964_ = ~new_n1963_;
  assign new_n1965_ = new_n951_ & new_n279_;
  assign new_n1966_ = ~new_n1965_;
  assign new_n1967_ = new_n1966_ & new_n1964_;
  assign new_n1968_ = new_n1967_ & new_n318_;
  assign new_n1969_ = ~new_n1968_;
  assign new_n1970_ = new_n961_ & shift1;
  assign new_n1971_ = ~new_n1970_;
  assign new_n1972_ = new_n904_ & new_n279_;
  assign new_n1973_ = ~new_n1972_;
  assign new_n1974_ = new_n1973_ & new_n1971_;
  assign new_n1975_ = new_n1974_ & new_n342_;
  assign new_n1976_ = ~new_n1975_;
  assign new_n1977_ = new_n1976_ & new_n1969_;
  assign new_n1978_ = new_n1977_ & new_n1962_;
  assign new_n1979_ = ~new_n1978_;
  assign new_n1980_ = new_n1979_ & new_n570_;
  assign new_n1981_ = ~new_n1980_;
  assign new_n1982_ = new_n694_ & shift1;
  assign new_n1983_ = ~new_n1982_;
  assign new_n1984_ = new_n829_ & new_n279_;
  assign new_n1985_ = ~new_n1984_;
  assign new_n1986_ = new_n1985_ & new_n1983_;
  assign new_n1987_ = new_n1986_ & new_n267_;
  assign new_n1988_ = ~new_n1987_;
  assign new_n1989_ = new_n717_ & shift1;
  assign new_n1990_ = ~new_n1989_;
  assign new_n1991_ = new_n684_ & new_n279_;
  assign new_n1992_ = ~new_n1991_;
  assign new_n1993_ = new_n1992_ & new_n1990_;
  assign new_n1994_ = new_n1993_ & new_n293_;
  assign new_n1995_ = ~new_n1994_;
  assign new_n1996_ = new_n1995_ & new_n1988_;
  assign new_n1997_ = new_n741_ & shift1;
  assign new_n1998_ = ~new_n1997_;
  assign new_n1999_ = new_n754_ & new_n279_;
  assign new_n2000_ = ~new_n1999_;
  assign new_n2001_ = new_n2000_ & new_n1998_;
  assign new_n2002_ = new_n2001_ & new_n318_;
  assign new_n2003_ = ~new_n2002_;
  assign new_n2004_ = new_n764_ & shift1;
  assign new_n2005_ = ~new_n2004_;
  assign new_n2006_ = new_n707_ & new_n279_;
  assign new_n2007_ = ~new_n2006_;
  assign new_n2008_ = new_n2007_ & new_n2005_;
  assign new_n2009_ = new_n2008_ & new_n342_;
  assign new_n2010_ = ~new_n2009_;
  assign new_n2011_ = new_n2010_ & new_n2003_;
  assign new_n2012_ = new_n2011_ & new_n1996_;
  assign new_n2013_ = ~new_n2012_;
  assign new_n2014_ = new_n2013_ & new_n369_;
  assign new_n2015_ = ~new_n2014_;
  assign new_n2016_ = new_n2015_ & new_n1981_;
  assign new_n2017_ = new_n989_ & shift1;
  assign new_n2018_ = ~new_n2017_;
  assign new_n2019_ = new_n928_ & new_n279_;
  assign new_n2020_ = ~new_n2019_;
  assign new_n2021_ = new_n2020_ & new_n2018_;
  assign new_n2022_ = new_n2021_ & new_n267_;
  assign new_n2023_ = ~new_n2022_;
  assign new_n2024_ = new_n1012_ & shift1;
  assign new_n2025_ = ~new_n2024_;
  assign new_n2026_ = new_n979_ & new_n279_;
  assign new_n2027_ = ~new_n2026_;
  assign new_n2028_ = new_n2027_ & new_n2025_;
  assign new_n2029_ = new_n2028_ & new_n293_;
  assign new_n2030_ = ~new_n2029_;
  assign new_n2031_ = new_n2030_ & new_n2023_;
  assign new_n2032_ = ~new_n1052_;
  assign new_n2033_ = new_n2032_ & new_n1047_;
  assign new_n2034_ = ~new_n2033_;
  assign new_n2035_ = new_n2034_ & new_n279_;
  assign new_n2036_ = ~new_n2035_;
  assign new_n2037_ = new_n1035_ & shift1;
  assign new_n2038_ = ~new_n2037_;
  assign new_n2039_ = new_n2038_ & new_n2036_;
  assign new_n2040_ = ~new_n2039_;
  assign new_n2041_ = new_n2040_ & new_n318_;
  assign new_n2042_ = ~new_n2041_;
  assign new_n2043_ = new_n1001_ & new_n279_;
  assign new_n2044_ = ~new_n2043_;
  assign new_n2045_ = ~new_n1055_;
  assign new_n2046_ = new_n2045_ & new_n1043_;
  assign new_n2047_ = ~new_n2046_;
  assign new_n2048_ = new_n2047_ & shift1;
  assign new_n2049_ = ~new_n2048_;
  assign new_n2050_ = new_n2049_ & new_n2044_;
  assign new_n2051_ = ~new_n2050_;
  assign new_n2052_ = new_n2051_ & new_n342_;
  assign new_n2053_ = ~new_n2052_;
  assign new_n2054_ = new_n2053_ & new_n2042_;
  assign new_n2055_ = new_n2054_ & new_n2031_;
  assign new_n2056_ = ~new_n2055_;
  assign new_n2057_ = new_n2056_ & new_n669_;
  assign new_n2058_ = ~new_n2057_;
  assign new_n2059_ = new_n792_ & shift1;
  assign new_n2060_ = ~new_n2059_;
  assign new_n2061_ = new_n1026_ & new_n279_;
  assign new_n2062_ = ~new_n2061_;
  assign new_n2063_ = new_n2062_ & new_n2060_;
  assign new_n2064_ = new_n2063_ & new_n267_;
  assign new_n2065_ = ~new_n2064_;
  assign new_n2066_ = new_n815_ & shift1;
  assign new_n2067_ = ~new_n2066_;
  assign new_n2068_ = new_n782_ & new_n279_;
  assign new_n2069_ = ~new_n2068_;
  assign new_n2070_ = new_n2069_ & new_n2067_;
  assign new_n2071_ = new_n2070_ & new_n293_;
  assign new_n2072_ = ~new_n2071_;
  assign new_n2073_ = new_n2072_ & new_n2065_;
  assign new_n2074_ = new_n839_ & shift1;
  assign new_n2075_ = ~new_n2074_;
  assign new_n2076_ = new_n852_ & new_n279_;
  assign new_n2077_ = ~new_n2076_;
  assign new_n2078_ = new_n2077_ & new_n2075_;
  assign new_n2079_ = new_n2078_ & new_n318_;
  assign new_n2080_ = ~new_n2079_;
  assign new_n2081_ = new_n862_ & shift1;
  assign new_n2082_ = ~new_n2081_;
  assign new_n2083_ = new_n805_ & new_n279_;
  assign new_n2084_ = ~new_n2083_;
  assign new_n2085_ = new_n2084_ & new_n2082_;
  assign new_n2086_ = new_n2085_ & new_n342_;
  assign new_n2087_ = ~new_n2086_;
  assign new_n2088_ = new_n2087_ & new_n2080_;
  assign new_n2089_ = new_n2088_ & new_n2073_;
  assign new_n2090_ = ~new_n2089_;
  assign new_n2091_ = new_n2090_ & new_n469_;
  assign new_n2092_ = ~new_n2091_;
  assign new_n2093_ = new_n2092_ & new_n2058_;
  assign new_n2094_ = new_n2093_ & new_n2016_;
  assign new_n2095_ = ~new_n2094_;
  assign new_n2096_ = new_n2095_ & shift6;
  assign new_n2097_ = ~new_n2096_;
  assign new_n2098_ = new_n2097_ & new_n1947_;
  assign ores2 = ~new_n2098_;
  assign new_n2100_ = new_n1304_ & new_n279_;
  assign new_n2101_ = ~new_n2100_;
  assign new_n2102_ = new_n1347_ & shift1;
  assign new_n2103_ = ~new_n2102_;
  assign new_n2104_ = new_n2103_ & new_n2101_;
  assign new_n2105_ = ~new_n2104_;
  assign new_n2106_ = new_n1359_ & shift1;
  assign new_n2107_ = ~new_n2106_;
  assign new_n2108_ = new_n1309_ & new_n279_;
  assign new_n2109_ = ~new_n2108_;
  assign new_n2110_ = new_n2109_ & new_n2107_;
  assign new_n2111_ = new_n2110_ & new_n2105_;
  assign new_n2112_ = ~new_n2111_;
  assign new_n2113_ = new_n2112_ & new_n267_;
  assign new_n2114_ = ~new_n2113_;
  assign new_n2115_ = new_n1351_ & new_n279_;
  assign new_n2116_ = ~new_n2115_;
  assign new_n2117_ = new_n1368_ & shift1;
  assign new_n2118_ = ~new_n2117_;
  assign new_n2119_ = new_n2118_ & new_n2116_;
  assign new_n2120_ = ~new_n2119_;
  assign new_n2121_ = new_n1380_ & shift1;
  assign new_n2122_ = ~new_n2121_;
  assign new_n2123_ = new_n1356_ & new_n279_;
  assign new_n2124_ = ~new_n2123_;
  assign new_n2125_ = new_n2124_ & new_n2122_;
  assign new_n2126_ = new_n2125_ & new_n2120_;
  assign new_n2127_ = ~new_n2126_;
  assign new_n2128_ = new_n2127_ & new_n293_;
  assign new_n2129_ = ~new_n2128_;
  assign new_n2130_ = new_n2129_ & new_n2114_;
  assign new_n2131_ = new_n1415_ & new_n279_;
  assign new_n2132_ = ~new_n2131_;
  assign new_n2133_ = new_n1390_ & shift1;
  assign new_n2134_ = ~new_n2133_;
  assign new_n2135_ = new_n2134_ & new_n2132_;
  assign new_n2136_ = ~new_n2135_;
  assign new_n2137_ = new_n1402_ & shift1;
  assign new_n2138_ = ~new_n2137_;
  assign new_n2139_ = new_n1420_ & new_n279_;
  assign new_n2140_ = ~new_n2139_;
  assign new_n2141_ = new_n2140_ & new_n2138_;
  assign new_n2142_ = new_n2141_ & new_n2136_;
  assign new_n2143_ = ~new_n2142_;
  assign new_n2144_ = new_n2143_ & new_n318_;
  assign new_n2145_ = ~new_n2144_;
  assign new_n2146_ = new_n1372_ & new_n279_;
  assign new_n2147_ = ~new_n2146_;
  assign new_n2148_ = new_n1411_ & shift1;
  assign new_n2149_ = ~new_n2148_;
  assign new_n2150_ = new_n2149_ & new_n2147_;
  assign new_n2151_ = ~new_n2150_;
  assign new_n2152_ = new_n1423_ & shift1;
  assign new_n2153_ = ~new_n2152_;
  assign new_n2154_ = new_n1377_ & new_n279_;
  assign new_n2155_ = ~new_n2154_;
  assign new_n2156_ = new_n2155_ & new_n2153_;
  assign new_n2157_ = new_n2156_ & new_n2151_;
  assign new_n2158_ = ~new_n2157_;
  assign new_n2159_ = new_n2158_ & new_n342_;
  assign new_n2160_ = ~new_n2159_;
  assign new_n2161_ = new_n2160_ & new_n2145_;
  assign new_n2162_ = new_n2161_ & new_n2130_;
  assign new_n2163_ = ~new_n2162_;
  assign new_n2164_ = new_n2163_ & new_n669_;
  assign new_n2165_ = ~new_n2164_;
  assign new_n2166_ = new_n1394_ & new_n279_;
  assign new_n2167_ = ~new_n2166_;
  assign new_n2168_ = new_n1166_ & shift1;
  assign new_n2169_ = ~new_n2168_;
  assign new_n2170_ = new_n2169_ & new_n2167_;
  assign new_n2171_ = ~new_n2170_;
  assign new_n2172_ = new_n1178_ & shift1;
  assign new_n2173_ = ~new_n2172_;
  assign new_n2174_ = new_n1399_ & new_n279_;
  assign new_n2175_ = ~new_n2174_;
  assign new_n2176_ = new_n2175_ & new_n2173_;
  assign new_n2177_ = new_n2176_ & new_n2171_;
  assign new_n2178_ = ~new_n2177_;
  assign new_n2179_ = new_n2178_ & new_n267_;
  assign new_n2180_ = ~new_n2179_;
  assign new_n2181_ = new_n1170_ & new_n279_;
  assign new_n2182_ = ~new_n2181_;
  assign new_n2183_ = new_n1187_ & shift1;
  assign new_n2184_ = ~new_n2183_;
  assign new_n2185_ = new_n2184_ & new_n2182_;
  assign new_n2186_ = ~new_n2185_;
  assign new_n2187_ = new_n1199_ & shift1;
  assign new_n2188_ = ~new_n2187_;
  assign new_n2189_ = new_n1175_ & new_n279_;
  assign new_n2190_ = ~new_n2189_;
  assign new_n2191_ = new_n2190_ & new_n2188_;
  assign new_n2192_ = new_n2191_ & new_n2186_;
  assign new_n2193_ = ~new_n2192_;
  assign new_n2194_ = new_n2193_ & new_n293_;
  assign new_n2195_ = ~new_n2194_;
  assign new_n2196_ = new_n2195_ & new_n2180_;
  assign new_n2197_ = new_n1234_ & new_n279_;
  assign new_n2198_ = ~new_n2197_;
  assign new_n2199_ = new_n1209_ & shift1;
  assign new_n2200_ = ~new_n2199_;
  assign new_n2201_ = new_n2200_ & new_n2198_;
  assign new_n2202_ = ~new_n2201_;
  assign new_n2203_ = new_n1221_ & shift1;
  assign new_n2204_ = ~new_n2203_;
  assign new_n2205_ = new_n1239_ & new_n279_;
  assign new_n2206_ = ~new_n2205_;
  assign new_n2207_ = new_n2206_ & new_n2204_;
  assign new_n2208_ = new_n2207_ & new_n2202_;
  assign new_n2209_ = ~new_n2208_;
  assign new_n2210_ = new_n2209_ & new_n318_;
  assign new_n2211_ = ~new_n2210_;
  assign new_n2212_ = new_n1191_ & new_n279_;
  assign new_n2213_ = ~new_n2212_;
  assign new_n2214_ = new_n1230_ & shift1;
  assign new_n2215_ = ~new_n2214_;
  assign new_n2216_ = new_n2215_ & new_n2213_;
  assign new_n2217_ = ~new_n2216_;
  assign new_n2218_ = new_n1242_ & shift1;
  assign new_n2219_ = ~new_n2218_;
  assign new_n2220_ = new_n1196_ & new_n279_;
  assign new_n2221_ = ~new_n2220_;
  assign new_n2222_ = new_n2221_ & new_n2219_;
  assign new_n2223_ = new_n2222_ & new_n2217_;
  assign new_n2224_ = ~new_n2223_;
  assign new_n2225_ = new_n2224_ & new_n342_;
  assign new_n2226_ = ~new_n2225_;
  assign new_n2227_ = new_n2226_ & new_n2211_;
  assign new_n2228_ = new_n2227_ & new_n2196_;
  assign new_n2229_ = ~new_n2228_;
  assign new_n2230_ = new_n2229_ & new_n469_;
  assign new_n2231_ = ~new_n2230_;
  assign new_n2232_ = new_n2231_ & new_n2165_;
  assign new_n2233_ = new_n1579_ & new_n279_;
  assign new_n2234_ = ~new_n2233_;
  assign new_n2235_ = new_n1257_ & shift1;
  assign new_n2236_ = ~new_n2235_;
  assign new_n2237_ = new_n2236_ & new_n2234_;
  assign new_n2238_ = ~new_n2237_;
  assign new_n2239_ = new_n1269_ & shift1;
  assign new_n2240_ = ~new_n2239_;
  assign new_n2241_ = new_n1584_ & new_n279_;
  assign new_n2242_ = ~new_n2241_;
  assign new_n2243_ = new_n2242_ & new_n2240_;
  assign new_n2244_ = new_n2243_ & new_n2238_;
  assign new_n2245_ = ~new_n2244_;
  assign new_n2246_ = new_n2245_ & new_n267_;
  assign new_n2247_ = ~new_n2246_;
  assign new_n2248_ = new_n1261_ & new_n279_;
  assign new_n2249_ = ~new_n2248_;
  assign new_n2250_ = new_n1278_ & shift1;
  assign new_n2251_ = ~new_n2250_;
  assign new_n2252_ = new_n2251_ & new_n2249_;
  assign new_n2253_ = ~new_n2252_;
  assign new_n2254_ = new_n1290_ & shift1;
  assign new_n2255_ = ~new_n2254_;
  assign new_n2256_ = new_n1266_ & new_n279_;
  assign new_n2257_ = ~new_n2256_;
  assign new_n2258_ = new_n2257_ & new_n2255_;
  assign new_n2259_ = new_n2258_ & new_n2253_;
  assign new_n2260_ = ~new_n2259_;
  assign new_n2261_ = new_n2260_ & new_n293_;
  assign new_n2262_ = ~new_n2261_;
  assign new_n2263_ = new_n2262_ & new_n2247_;
  assign new_n2264_ = new_n1325_ & new_n279_;
  assign new_n2265_ = ~new_n2264_;
  assign new_n2266_ = new_n1300_ & shift1;
  assign new_n2267_ = ~new_n2266_;
  assign new_n2268_ = new_n2267_ & new_n2265_;
  assign new_n2269_ = ~new_n2268_;
  assign new_n2270_ = new_n1312_ & shift1;
  assign new_n2271_ = ~new_n2270_;
  assign new_n2272_ = new_n1330_ & new_n279_;
  assign new_n2273_ = ~new_n2272_;
  assign new_n2274_ = new_n2273_ & new_n2271_;
  assign new_n2275_ = new_n2274_ & new_n2269_;
  assign new_n2276_ = ~new_n2275_;
  assign new_n2277_ = new_n2276_ & new_n318_;
  assign new_n2278_ = ~new_n2277_;
  assign new_n2279_ = new_n1282_ & new_n279_;
  assign new_n2280_ = ~new_n2279_;
  assign new_n2281_ = new_n1321_ & shift1;
  assign new_n2282_ = ~new_n2281_;
  assign new_n2283_ = new_n2282_ & new_n2280_;
  assign new_n2284_ = ~new_n2283_;
  assign new_n2285_ = new_n1333_ & shift1;
  assign new_n2286_ = ~new_n2285_;
  assign new_n2287_ = new_n1287_ & new_n279_;
  assign new_n2288_ = ~new_n2287_;
  assign new_n2289_ = new_n2288_ & new_n2286_;
  assign new_n2290_ = new_n2289_ & new_n2284_;
  assign new_n2291_ = ~new_n2290_;
  assign new_n2292_ = new_n2291_ & new_n342_;
  assign new_n2293_ = ~new_n2292_;
  assign new_n2294_ = new_n2293_ & new_n2278_;
  assign new_n2295_ = new_n2294_ & new_n2263_;
  assign new_n2296_ = ~new_n2295_;
  assign new_n2297_ = new_n2296_ & new_n570_;
  assign new_n2298_ = ~new_n2297_;
  assign new_n2299_ = new_n1213_ & new_n279_;
  assign new_n2300_ = ~new_n2299_;
  assign new_n2301_ = new_n1076_ & shift1;
  assign new_n2302_ = ~new_n2301_;
  assign new_n2303_ = new_n2302_ & new_n2300_;
  assign new_n2304_ = ~new_n2303_;
  assign new_n2305_ = new_n1088_ & shift1;
  assign new_n2306_ = ~new_n2305_;
  assign new_n2307_ = new_n1218_ & new_n279_;
  assign new_n2308_ = ~new_n2307_;
  assign new_n2309_ = new_n2308_ & new_n2306_;
  assign new_n2310_ = new_n2309_ & new_n2304_;
  assign new_n2311_ = ~new_n2310_;
  assign new_n2312_ = new_n2311_ & new_n267_;
  assign new_n2313_ = ~new_n2312_;
  assign new_n2314_ = new_n1080_ & new_n279_;
  assign new_n2315_ = ~new_n2314_;
  assign new_n2316_ = new_n1097_ & shift1;
  assign new_n2317_ = ~new_n2316_;
  assign new_n2318_ = new_n2317_ & new_n2315_;
  assign new_n2319_ = ~new_n2318_;
  assign new_n2320_ = new_n1109_ & shift1;
  assign new_n2321_ = ~new_n2320_;
  assign new_n2322_ = new_n1085_ & new_n279_;
  assign new_n2323_ = ~new_n2322_;
  assign new_n2324_ = new_n2323_ & new_n2321_;
  assign new_n2325_ = new_n2324_ & new_n2319_;
  assign new_n2326_ = ~new_n2325_;
  assign new_n2327_ = new_n2326_ & new_n293_;
  assign new_n2328_ = ~new_n2327_;
  assign new_n2329_ = new_n2328_ & new_n2313_;
  assign new_n2330_ = new_n1144_ & new_n279_;
  assign new_n2331_ = ~new_n2330_;
  assign new_n2332_ = new_n1119_ & shift1;
  assign new_n2333_ = ~new_n2332_;
  assign new_n2334_ = new_n2333_ & new_n2331_;
  assign new_n2335_ = ~new_n2334_;
  assign new_n2336_ = new_n1131_ & shift1;
  assign new_n2337_ = ~new_n2336_;
  assign new_n2338_ = new_n1149_ & new_n279_;
  assign new_n2339_ = ~new_n2338_;
  assign new_n2340_ = new_n2339_ & new_n2337_;
  assign new_n2341_ = new_n2340_ & new_n2335_;
  assign new_n2342_ = ~new_n2341_;
  assign new_n2343_ = new_n2342_ & new_n318_;
  assign new_n2344_ = ~new_n2343_;
  assign new_n2345_ = new_n1101_ & new_n279_;
  assign new_n2346_ = ~new_n2345_;
  assign new_n2347_ = new_n1140_ & shift1;
  assign new_n2348_ = ~new_n2347_;
  assign new_n2349_ = new_n2348_ & new_n2346_;
  assign new_n2350_ = ~new_n2349_;
  assign new_n2351_ = new_n1152_ & shift1;
  assign new_n2352_ = ~new_n2351_;
  assign new_n2353_ = new_n1106_ & new_n279_;
  assign new_n2354_ = ~new_n2353_;
  assign new_n2355_ = new_n2354_ & new_n2352_;
  assign new_n2356_ = new_n2355_ & new_n2350_;
  assign new_n2357_ = ~new_n2356_;
  assign new_n2358_ = new_n2357_ & new_n342_;
  assign new_n2359_ = ~new_n2358_;
  assign new_n2360_ = new_n2359_ & new_n2344_;
  assign new_n2361_ = new_n2360_ & new_n2329_;
  assign new_n2362_ = ~new_n2361_;
  assign new_n2363_ = new_n2362_ & new_n369_;
  assign new_n2364_ = ~new_n2363_;
  assign new_n2365_ = new_n2364_ & new_n2298_;
  assign new_n2366_ = new_n2365_ & new_n2232_;
  assign new_n2367_ = ~new_n2366_;
  assign new_n2368_ = new_n2367_ & new_n264_;
  assign new_n2369_ = ~new_n2368_;
  assign new_n2370_ = new_n1123_ & new_n279_;
  assign new_n2371_ = ~new_n2370_;
  assign new_n2372_ = new_n1442_ & shift1;
  assign new_n2373_ = ~new_n2372_;
  assign new_n2374_ = new_n2373_ & new_n2371_;
  assign new_n2375_ = ~new_n2374_;
  assign new_n2376_ = new_n1454_ & shift1;
  assign new_n2377_ = ~new_n2376_;
  assign new_n2378_ = new_n1128_ & new_n279_;
  assign new_n2379_ = ~new_n2378_;
  assign new_n2380_ = new_n2379_ & new_n2377_;
  assign new_n2381_ = new_n2380_ & new_n2375_;
  assign new_n2382_ = ~new_n2381_;
  assign new_n2383_ = new_n2382_ & new_n267_;
  assign new_n2384_ = ~new_n2383_;
  assign new_n2385_ = new_n1446_ & new_n279_;
  assign new_n2386_ = ~new_n2385_;
  assign new_n2387_ = new_n1463_ & shift1;
  assign new_n2388_ = ~new_n2387_;
  assign new_n2389_ = new_n2388_ & new_n2386_;
  assign new_n2390_ = ~new_n2389_;
  assign new_n2391_ = new_n1475_ & shift1;
  assign new_n2392_ = ~new_n2391_;
  assign new_n2393_ = new_n1451_ & new_n279_;
  assign new_n2394_ = ~new_n2393_;
  assign new_n2395_ = new_n2394_ & new_n2392_;
  assign new_n2396_ = new_n2395_ & new_n2390_;
  assign new_n2397_ = ~new_n2396_;
  assign new_n2398_ = new_n2397_ & new_n293_;
  assign new_n2399_ = ~new_n2398_;
  assign new_n2400_ = new_n2399_ & new_n2384_;
  assign new_n2401_ = new_n1510_ & new_n279_;
  assign new_n2402_ = ~new_n2401_;
  assign new_n2403_ = new_n1485_ & shift1;
  assign new_n2404_ = ~new_n2403_;
  assign new_n2405_ = new_n2404_ & new_n2402_;
  assign new_n2406_ = ~new_n2405_;
  assign new_n2407_ = new_n1497_ & shift1;
  assign new_n2408_ = ~new_n2407_;
  assign new_n2409_ = new_n1515_ & new_n279_;
  assign new_n2410_ = ~new_n2409_;
  assign new_n2411_ = new_n2410_ & new_n2408_;
  assign new_n2412_ = new_n2411_ & new_n2406_;
  assign new_n2413_ = ~new_n2412_;
  assign new_n2414_ = new_n2413_ & new_n318_;
  assign new_n2415_ = ~new_n2414_;
  assign new_n2416_ = new_n1467_ & new_n279_;
  assign new_n2417_ = ~new_n2416_;
  assign new_n2418_ = new_n1506_ & shift1;
  assign new_n2419_ = ~new_n2418_;
  assign new_n2420_ = new_n2419_ & new_n2417_;
  assign new_n2421_ = ~new_n2420_;
  assign new_n2422_ = new_n1518_ & shift1;
  assign new_n2423_ = ~new_n2422_;
  assign new_n2424_ = new_n1472_ & new_n279_;
  assign new_n2425_ = ~new_n2424_;
  assign new_n2426_ = new_n2425_ & new_n2423_;
  assign new_n2427_ = new_n2426_ & new_n2421_;
  assign new_n2428_ = ~new_n2427_;
  assign new_n2429_ = new_n2428_ & new_n342_;
  assign new_n2430_ = ~new_n2429_;
  assign new_n2431_ = new_n2430_ & new_n2415_;
  assign new_n2432_ = new_n2431_ & new_n2400_;
  assign new_n2433_ = ~new_n2432_;
  assign new_n2434_ = new_n2433_ & new_n570_;
  assign new_n2435_ = ~new_n2434_;
  assign new_n2436_ = new_n1489_ & new_n279_;
  assign new_n2437_ = ~new_n2436_;
  assign new_n2438_ = new_n1623_ & shift1;
  assign new_n2439_ = ~new_n2438_;
  assign new_n2440_ = new_n2439_ & new_n2437_;
  assign new_n2441_ = ~new_n2440_;
  assign new_n2442_ = new_n1635_ & shift1;
  assign new_n2443_ = ~new_n2442_;
  assign new_n2444_ = new_n1494_ & new_n279_;
  assign new_n2445_ = ~new_n2444_;
  assign new_n2446_ = new_n2445_ & new_n2443_;
  assign new_n2447_ = new_n2446_ & new_n2441_;
  assign new_n2448_ = ~new_n2447_;
  assign new_n2449_ = new_n2448_ & new_n267_;
  assign new_n2450_ = ~new_n2449_;
  assign new_n2451_ = new_n1655_ & shift1;
  assign new_n2452_ = ~new_n2451_;
  assign new_n2453_ = ~new_n1632_;
  assign new_n2454_ = new_n2453_ & new_n1627_;
  assign new_n2455_ = ~new_n2454_;
  assign new_n2456_ = new_n2455_ & new_n279_;
  assign new_n2457_ = ~new_n2456_;
  assign new_n2458_ = new_n2457_ & new_n2452_;
  assign new_n2459_ = ~new_n2458_;
  assign new_n2460_ = new_n2459_ & new_n293_;
  assign new_n2461_ = ~new_n2460_;
  assign new_n2462_ = new_n2461_ & new_n2450_;
  assign new_n2463_ = new_n1693_ & new_n279_;
  assign new_n2464_ = ~new_n2463_;
  assign new_n2465_ = new_n1664_ & shift1;
  assign new_n2466_ = ~new_n2465_;
  assign new_n2467_ = new_n2466_ & new_n2464_;
  assign new_n2468_ = ~new_n2467_;
  assign new_n2469_ = new_n1676_ & shift1;
  assign new_n2470_ = ~new_n2469_;
  assign new_n2471_ = new_n1694_ & new_n279_;
  assign new_n2472_ = ~new_n2471_;
  assign new_n2473_ = new_n2472_ & new_n2470_;
  assign new_n2474_ = new_n2473_ & new_n2468_;
  assign new_n2475_ = ~new_n2474_;
  assign new_n2476_ = new_n2475_ & new_n318_;
  assign new_n2477_ = ~new_n2476_;
  assign new_n2478_ = new_n1646_ & new_n279_;
  assign new_n2479_ = ~new_n2478_;
  assign new_n2480_ = new_n1687_ & shift1;
  assign new_n2481_ = ~new_n2480_;
  assign new_n2482_ = new_n2481_ & new_n2479_;
  assign new_n2483_ = ~new_n2482_;
  assign new_n2484_ = new_n1684_ & shift1;
  assign new_n2485_ = ~new_n2484_;
  assign new_n2486_ = new_n1643_ & new_n279_;
  assign new_n2487_ = ~new_n2486_;
  assign new_n2488_ = new_n2487_ & new_n2485_;
  assign new_n2489_ = new_n2488_ & new_n2483_;
  assign new_n2490_ = ~new_n2489_;
  assign new_n2491_ = new_n2490_ & new_n342_;
  assign new_n2492_ = ~new_n2491_;
  assign new_n2493_ = new_n2492_ & new_n2477_;
  assign new_n2494_ = new_n2493_ & new_n2462_;
  assign new_n2495_ = ~new_n2494_;
  assign new_n2496_ = new_n2495_ & new_n669_;
  assign new_n2497_ = ~new_n2496_;
  assign new_n2498_ = new_n2497_ & new_n2435_;
  assign new_n2499_ = new_n1757_ & new_n279_;
  assign new_n2500_ = ~new_n2499_;
  assign new_n2501_ = new_n1532_ & shift1;
  assign new_n2502_ = ~new_n2501_;
  assign new_n2503_ = new_n2502_ & new_n2500_;
  assign new_n2504_ = ~new_n2503_;
  assign new_n2505_ = new_n1544_ & shift1;
  assign new_n2506_ = ~new_n2505_;
  assign new_n2507_ = new_n1762_ & new_n279_;
  assign new_n2508_ = ~new_n2507_;
  assign new_n2509_ = new_n2508_ & new_n2506_;
  assign new_n2510_ = new_n2509_ & new_n2504_;
  assign new_n2511_ = ~new_n2510_;
  assign new_n2512_ = new_n2511_ & new_n267_;
  assign new_n2513_ = ~new_n2512_;
  assign new_n2514_ = new_n1536_ & new_n279_;
  assign new_n2515_ = ~new_n2514_;
  assign new_n2516_ = new_n1553_ & shift1;
  assign new_n2517_ = ~new_n2516_;
  assign new_n2518_ = new_n2517_ & new_n2515_;
  assign new_n2519_ = ~new_n2518_;
  assign new_n2520_ = new_n1565_ & shift1;
  assign new_n2521_ = ~new_n2520_;
  assign new_n2522_ = new_n1541_ & new_n279_;
  assign new_n2523_ = ~new_n2522_;
  assign new_n2524_ = new_n2523_ & new_n2521_;
  assign new_n2525_ = new_n2524_ & new_n2519_;
  assign new_n2526_ = ~new_n2525_;
  assign new_n2527_ = new_n2526_ & new_n293_;
  assign new_n2528_ = ~new_n2527_;
  assign new_n2529_ = new_n2528_ & new_n2513_;
  assign new_n2530_ = new_n1600_ & new_n279_;
  assign new_n2531_ = ~new_n2530_;
  assign new_n2532_ = new_n1575_ & shift1;
  assign new_n2533_ = ~new_n2532_;
  assign new_n2534_ = new_n2533_ & new_n2531_;
  assign new_n2535_ = ~new_n2534_;
  assign new_n2536_ = new_n1587_ & shift1;
  assign new_n2537_ = ~new_n2536_;
  assign new_n2538_ = new_n1605_ & new_n279_;
  assign new_n2539_ = ~new_n2538_;
  assign new_n2540_ = new_n2539_ & new_n2537_;
  assign new_n2541_ = new_n2540_ & new_n2535_;
  assign new_n2542_ = ~new_n2541_;
  assign new_n2543_ = new_n2542_ & new_n318_;
  assign new_n2544_ = ~new_n2543_;
  assign new_n2545_ = new_n1557_ & new_n279_;
  assign new_n2546_ = ~new_n2545_;
  assign new_n2547_ = new_n1596_ & shift1;
  assign new_n2548_ = ~new_n2547_;
  assign new_n2549_ = new_n2548_ & new_n2546_;
  assign new_n2550_ = ~new_n2549_;
  assign new_n2551_ = new_n1608_ & shift1;
  assign new_n2552_ = ~new_n2551_;
  assign new_n2553_ = new_n1562_ & new_n279_;
  assign new_n2554_ = ~new_n2553_;
  assign new_n2555_ = new_n2554_ & new_n2552_;
  assign new_n2556_ = new_n2555_ & new_n2550_;
  assign new_n2557_ = ~new_n2556_;
  assign new_n2558_ = new_n2557_ & new_n342_;
  assign new_n2559_ = ~new_n2558_;
  assign new_n2560_ = new_n2559_ & new_n2544_;
  assign new_n2561_ = new_n2560_ & new_n2529_;
  assign new_n2562_ = ~new_n2561_;
  assign new_n2563_ = new_n2562_ & new_n369_;
  assign new_n2564_ = ~new_n2563_;
  assign new_n2565_ = new_n1668_ & new_n279_;
  assign new_n2566_ = ~new_n2565_;
  assign new_n2567_ = new_n1710_ & shift1;
  assign new_n2568_ = ~new_n2567_;
  assign new_n2569_ = new_n2568_ & new_n2566_;
  assign new_n2570_ = ~new_n2569_;
  assign new_n2571_ = new_n1722_ & shift1;
  assign new_n2572_ = ~new_n2571_;
  assign new_n2573_ = new_n1673_ & new_n279_;
  assign new_n2574_ = ~new_n2573_;
  assign new_n2575_ = new_n2574_ & new_n2572_;
  assign new_n2576_ = new_n2575_ & new_n2570_;
  assign new_n2577_ = ~new_n2576_;
  assign new_n2578_ = new_n2577_ & new_n267_;
  assign new_n2579_ = ~new_n2578_;
  assign new_n2580_ = new_n1714_ & new_n279_;
  assign new_n2581_ = ~new_n2580_;
  assign new_n2582_ = new_n1731_ & shift1;
  assign new_n2583_ = ~new_n2582_;
  assign new_n2584_ = new_n2583_ & new_n2581_;
  assign new_n2585_ = ~new_n2584_;
  assign new_n2586_ = new_n1743_ & shift1;
  assign new_n2587_ = ~new_n2586_;
  assign new_n2588_ = new_n1719_ & new_n279_;
  assign new_n2589_ = ~new_n2588_;
  assign new_n2590_ = new_n2589_ & new_n2587_;
  assign new_n2591_ = new_n2590_ & new_n2585_;
  assign new_n2592_ = ~new_n2591_;
  assign new_n2593_ = new_n2592_ & new_n293_;
  assign new_n2594_ = ~new_n2593_;
  assign new_n2595_ = new_n2594_ & new_n2579_;
  assign new_n2596_ = new_n1778_ & new_n279_;
  assign new_n2597_ = ~new_n2596_;
  assign new_n2598_ = new_n1753_ & shift1;
  assign new_n2599_ = ~new_n2598_;
  assign new_n2600_ = new_n2599_ & new_n2597_;
  assign new_n2601_ = ~new_n2600_;
  assign new_n2602_ = new_n1765_ & shift1;
  assign new_n2603_ = ~new_n2602_;
  assign new_n2604_ = new_n1783_ & new_n279_;
  assign new_n2605_ = ~new_n2604_;
  assign new_n2606_ = new_n2605_ & new_n2603_;
  assign new_n2607_ = new_n2606_ & new_n2601_;
  assign new_n2608_ = ~new_n2607_;
  assign new_n2609_ = new_n2608_ & new_n318_;
  assign new_n2610_ = ~new_n2609_;
  assign new_n2611_ = new_n1735_ & new_n279_;
  assign new_n2612_ = ~new_n2611_;
  assign new_n2613_ = new_n1774_ & shift1;
  assign new_n2614_ = ~new_n2613_;
  assign new_n2615_ = new_n2614_ & new_n2612_;
  assign new_n2616_ = ~new_n2615_;
  assign new_n2617_ = new_n1786_ & shift1;
  assign new_n2618_ = ~new_n2617_;
  assign new_n2619_ = new_n1740_ & new_n279_;
  assign new_n2620_ = ~new_n2619_;
  assign new_n2621_ = new_n2620_ & new_n2618_;
  assign new_n2622_ = new_n2621_ & new_n2616_;
  assign new_n2623_ = ~new_n2622_;
  assign new_n2624_ = new_n2623_ & new_n342_;
  assign new_n2625_ = ~new_n2624_;
  assign new_n2626_ = new_n2625_ & new_n2610_;
  assign new_n2627_ = new_n2626_ & new_n2595_;
  assign new_n2628_ = ~new_n2627_;
  assign new_n2629_ = new_n2628_ & new_n469_;
  assign new_n2630_ = ~new_n2629_;
  assign new_n2631_ = new_n2630_ & new_n2564_;
  assign new_n2632_ = new_n2631_ & new_n2498_;
  assign new_n2633_ = ~new_n2632_;
  assign new_n2634_ = new_n2633_ & shift6;
  assign new_n2635_ = ~new_n2634_;
  assign new_n2636_ = new_n2635_ & new_n2369_;
  assign ores3 = ~new_n2636_;
  assign new_n2638_ = new_n439_ & new_n267_;
  assign new_n2639_ = ~new_n2638_;
  assign new_n2640_ = new_n293_ & new_n290_;
  assign new_n2641_ = ~new_n2640_;
  assign new_n2642_ = new_n2641_ & new_n2639_;
  assign new_n2643_ = new_n363_ & new_n318_;
  assign new_n2644_ = ~new_n2643_;
  assign new_n2645_ = new_n342_ & new_n314_;
  assign new_n2646_ = ~new_n2645_;
  assign new_n2647_ = new_n2646_ & new_n2644_;
  assign new_n2648_ = new_n2647_ & new_n2642_;
  assign new_n2649_ = ~new_n2648_;
  assign new_n2650_ = new_n2649_ & new_n369_;
  assign new_n2651_ = ~new_n2650_;
  assign new_n2652_ = new_n640_ & new_n267_;
  assign new_n2653_ = ~new_n2652_;
  assign new_n2654_ = new_n392_ & new_n293_;
  assign new_n2655_ = ~new_n2654_;
  assign new_n2656_ = new_n2655_ & new_n2653_;
  assign new_n2657_ = new_n462_ & new_n318_;
  assign new_n2658_ = ~new_n2657_;
  assign new_n2659_ = new_n415_ & new_n342_;
  assign new_n2660_ = ~new_n2659_;
  assign new_n2661_ = new_n2660_ & new_n2658_;
  assign new_n2662_ = new_n2661_ & new_n2656_;
  assign new_n2663_ = ~new_n2662_;
  assign new_n2664_ = new_n2663_ & new_n469_;
  assign new_n2665_ = ~new_n2664_;
  assign new_n2666_ = new_n2665_ & new_n2651_;
  assign new_n2667_ = new_n744_ & new_n267_;
  assign new_n2668_ = ~new_n2667_;
  assign new_n2669_ = new_n493_ & new_n293_;
  assign new_n2670_ = ~new_n2669_;
  assign new_n2671_ = new_n2670_ & new_n2668_;
  assign new_n2672_ = new_n563_ & new_n318_;
  assign new_n2673_ = ~new_n2672_;
  assign new_n2674_ = new_n516_ & new_n342_;
  assign new_n2675_ = ~new_n2674_;
  assign new_n2676_ = new_n2675_ & new_n2673_;
  assign new_n2677_ = new_n2676_ & new_n2671_;
  assign new_n2678_ = ~new_n2677_;
  assign new_n2679_ = new_n2678_ & new_n570_;
  assign new_n2680_ = ~new_n2679_;
  assign new_n2681_ = new_n540_ & new_n267_;
  assign new_n2682_ = ~new_n2681_;
  assign new_n2683_ = new_n593_ & new_n293_;
  assign new_n2684_ = ~new_n2683_;
  assign new_n2685_ = new_n2684_ & new_n2682_;
  assign new_n2686_ = new_n663_ & new_n318_;
  assign new_n2687_ = ~new_n2686_;
  assign new_n2688_ = new_n616_ & new_n342_;
  assign new_n2689_ = ~new_n2688_;
  assign new_n2690_ = new_n2689_ & new_n2687_;
  assign new_n2691_ = new_n2690_ & new_n2685_;
  assign new_n2692_ = ~new_n2691_;
  assign new_n2693_ = new_n2692_ & new_n669_;
  assign new_n2694_ = ~new_n2693_;
  assign new_n2695_ = new_n2694_ & new_n2680_;
  assign new_n2696_ = new_n2695_ & new_n2666_;
  assign new_n2697_ = ~new_n2696_;
  assign new_n2698_ = new_n2697_ & new_n264_;
  assign new_n2699_ = ~new_n2698_;
  assign new_n2700_ = new_n941_ & new_n267_;
  assign new_n2701_ = ~new_n2700_;
  assign new_n2702_ = new_n992_ & new_n293_;
  assign new_n2703_ = ~new_n2702_;
  assign new_n2704_ = new_n2703_ & new_n2701_;
  assign new_n2705_ = new_n1060_ & new_n318_;
  assign new_n2706_ = ~new_n2705_;
  assign new_n2707_ = new_n1015_ & new_n342_;
  assign new_n2708_ = ~new_n2707_;
  assign new_n2709_ = new_n2708_ & new_n2706_;
  assign new_n2710_ = new_n2709_ & new_n2704_;
  assign new_n2711_ = ~new_n2710_;
  assign new_n2712_ = new_n2711_ & new_n669_;
  assign new_n2713_ = ~new_n2712_;
  assign new_n2714_ = new_n339_ & new_n267_;
  assign new_n2715_ = ~new_n2714_;
  assign new_n2716_ = new_n894_ & new_n293_;
  assign new_n2717_ = ~new_n2716_;
  assign new_n2718_ = new_n2717_ & new_n2715_;
  assign new_n2719_ = new_n964_ & new_n318_;
  assign new_n2720_ = ~new_n2719_;
  assign new_n2721_ = new_n917_ & new_n342_;
  assign new_n2722_ = ~new_n2721_;
  assign new_n2723_ = new_n2722_ & new_n2720_;
  assign new_n2724_ = new_n2723_ & new_n2718_;
  assign new_n2725_ = ~new_n2724_;
  assign new_n2726_ = new_n2725_ & new_n570_;
  assign new_n2727_ = ~new_n2726_;
  assign new_n2728_ = new_n2727_ & new_n2713_;
  assign new_n2729_ = new_n1039_ & new_n267_;
  assign new_n2730_ = ~new_n2729_;
  assign new_n2731_ = new_n795_ & new_n293_;
  assign new_n2732_ = ~new_n2731_;
  assign new_n2733_ = new_n2732_ & new_n2730_;
  assign new_n2734_ = new_n865_ & new_n318_;
  assign new_n2735_ = ~new_n2734_;
  assign new_n2736_ = new_n818_ & new_n342_;
  assign new_n2737_ = ~new_n2736_;
  assign new_n2738_ = new_n2737_ & new_n2735_;
  assign new_n2739_ = new_n2738_ & new_n2733_;
  assign new_n2740_ = ~new_n2739_;
  assign new_n2741_ = new_n2740_ & new_n469_;
  assign new_n2742_ = ~new_n2741_;
  assign new_n2743_ = new_n842_ & new_n267_;
  assign new_n2744_ = ~new_n2743_;
  assign new_n2745_ = new_n697_ & new_n293_;
  assign new_n2746_ = ~new_n2745_;
  assign new_n2747_ = new_n2746_ & new_n2744_;
  assign new_n2748_ = new_n767_ & new_n318_;
  assign new_n2749_ = ~new_n2748_;
  assign new_n2750_ = new_n720_ & new_n342_;
  assign new_n2751_ = ~new_n2750_;
  assign new_n2752_ = new_n2751_ & new_n2749_;
  assign new_n2753_ = new_n2752_ & new_n2747_;
  assign new_n2754_ = ~new_n2753_;
  assign new_n2755_ = new_n2754_ & new_n369_;
  assign new_n2756_ = ~new_n2755_;
  assign new_n2757_ = new_n2756_ & new_n2742_;
  assign new_n2758_ = new_n2757_ & new_n2728_;
  assign new_n2759_ = ~new_n2758_;
  assign new_n2760_ = new_n2759_ & shift6;
  assign new_n2761_ = ~new_n2760_;
  assign new_n2762_ = new_n2761_ & new_n2699_;
  assign ores4 = ~new_n2762_;
  assign new_n2764_ = new_n1226_ & new_n267_;
  assign new_n2765_ = ~new_n2764_;
  assign new_n2766_ = new_n1093_ & new_n293_;
  assign new_n2767_ = ~new_n2766_;
  assign new_n2768_ = new_n2767_ & new_n2765_;
  assign new_n2769_ = new_n1157_ & new_n318_;
  assign new_n2770_ = ~new_n2769_;
  assign new_n2771_ = new_n1114_ & new_n342_;
  assign new_n2772_ = ~new_n2771_;
  assign new_n2773_ = new_n2772_ & new_n2770_;
  assign new_n2774_ = new_n2773_ & new_n2768_;
  assign new_n2775_ = ~new_n2774_;
  assign new_n2776_ = new_n2775_ & new_n369_;
  assign new_n2777_ = ~new_n2776_;
  assign new_n2778_ = new_n1407_ & new_n267_;
  assign new_n2779_ = ~new_n2778_;
  assign new_n2780_ = new_n1183_ & new_n293_;
  assign new_n2781_ = ~new_n2780_;
  assign new_n2782_ = new_n2781_ & new_n2779_;
  assign new_n2783_ = new_n1247_ & new_n318_;
  assign new_n2784_ = ~new_n2783_;
  assign new_n2785_ = new_n1204_ & new_n342_;
  assign new_n2786_ = ~new_n2785_;
  assign new_n2787_ = new_n2786_ & new_n2784_;
  assign new_n2788_ = new_n2787_ & new_n2782_;
  assign new_n2789_ = ~new_n2788_;
  assign new_n2790_ = new_n2789_ & new_n469_;
  assign new_n2791_ = ~new_n2790_;
  assign new_n2792_ = new_n2791_ & new_n2777_;
  assign new_n2793_ = new_n1592_ & new_n267_;
  assign new_n2794_ = ~new_n2793_;
  assign new_n2795_ = new_n1274_ & new_n293_;
  assign new_n2796_ = ~new_n2795_;
  assign new_n2797_ = new_n2796_ & new_n2794_;
  assign new_n2798_ = new_n1338_ & new_n318_;
  assign new_n2799_ = ~new_n2798_;
  assign new_n2800_ = new_n1295_ & new_n342_;
  assign new_n2801_ = ~new_n2800_;
  assign new_n2802_ = new_n2801_ & new_n2799_;
  assign new_n2803_ = new_n2802_ & new_n2797_;
  assign new_n2804_ = ~new_n2803_;
  assign new_n2805_ = new_n2804_ & new_n570_;
  assign new_n2806_ = ~new_n2805_;
  assign new_n2807_ = new_n1317_ & new_n267_;
  assign new_n2808_ = ~new_n2807_;
  assign new_n2809_ = new_n1364_ & new_n293_;
  assign new_n2810_ = ~new_n2809_;
  assign new_n2811_ = new_n2810_ & new_n2808_;
  assign new_n2812_ = new_n1428_ & new_n318_;
  assign new_n2813_ = ~new_n2812_;
  assign new_n2814_ = new_n1385_ & new_n342_;
  assign new_n2815_ = ~new_n2814_;
  assign new_n2816_ = new_n2815_ & new_n2813_;
  assign new_n2817_ = new_n2816_ & new_n2811_;
  assign new_n2818_ = ~new_n2817_;
  assign new_n2819_ = new_n2818_ & new_n669_;
  assign new_n2820_ = ~new_n2819_;
  assign new_n2821_ = new_n2820_ & new_n2806_;
  assign new_n2822_ = new_n2821_ & new_n2792_;
  assign new_n2823_ = ~new_n2822_;
  assign new_n2824_ = new_n2823_ & new_n264_;
  assign new_n2825_ = ~new_n2824_;
  assign new_n2826_ = new_n1502_ & new_n267_;
  assign new_n2827_ = ~new_n2826_;
  assign new_n2828_ = new_n1640_ & new_n293_;
  assign new_n2829_ = ~new_n2828_;
  assign new_n2830_ = new_n2829_ & new_n2827_;
  assign new_n2831_ = new_n1701_ & new_n318_;
  assign new_n2832_ = ~new_n2831_;
  assign new_n2833_ = new_n1659_ & new_n342_;
  assign new_n2834_ = ~new_n2833_;
  assign new_n2835_ = new_n2834_ & new_n2832_;
  assign new_n2836_ = new_n2835_ & new_n2830_;
  assign new_n2837_ = ~new_n2836_;
  assign new_n2838_ = new_n2837_ & new_n669_;
  assign new_n2839_ = ~new_n2838_;
  assign new_n2840_ = new_n1136_ & new_n267_;
  assign new_n2841_ = ~new_n2840_;
  assign new_n2842_ = new_n1459_ & new_n293_;
  assign new_n2843_ = ~new_n2842_;
  assign new_n2844_ = new_n2843_ & new_n2841_;
  assign new_n2845_ = new_n1523_ & new_n318_;
  assign new_n2846_ = ~new_n2845_;
  assign new_n2847_ = new_n1480_ & new_n342_;
  assign new_n2848_ = ~new_n2847_;
  assign new_n2849_ = new_n2848_ & new_n2846_;
  assign new_n2850_ = new_n2849_ & new_n2844_;
  assign new_n2851_ = ~new_n2850_;
  assign new_n2852_ = new_n2851_ & new_n570_;
  assign new_n2853_ = ~new_n2852_;
  assign new_n2854_ = new_n2853_ & new_n2839_;
  assign new_n2855_ = new_n1681_ & new_n267_;
  assign new_n2856_ = ~new_n2855_;
  assign new_n2857_ = new_n1727_ & new_n293_;
  assign new_n2858_ = ~new_n2857_;
  assign new_n2859_ = new_n2858_ & new_n2856_;
  assign new_n2860_ = new_n1791_ & new_n318_;
  assign new_n2861_ = ~new_n2860_;
  assign new_n2862_ = new_n1748_ & new_n342_;
  assign new_n2863_ = ~new_n2862_;
  assign new_n2864_ = new_n2863_ & new_n2861_;
  assign new_n2865_ = new_n2864_ & new_n2859_;
  assign new_n2866_ = ~new_n2865_;
  assign new_n2867_ = new_n2866_ & new_n469_;
  assign new_n2868_ = ~new_n2867_;
  assign new_n2869_ = new_n1770_ & new_n267_;
  assign new_n2870_ = ~new_n2869_;
  assign new_n2871_ = new_n1549_ & new_n293_;
  assign new_n2872_ = ~new_n2871_;
  assign new_n2873_ = new_n2872_ & new_n2870_;
  assign new_n2874_ = new_n1613_ & new_n318_;
  assign new_n2875_ = ~new_n2874_;
  assign new_n2876_ = new_n1570_ & new_n342_;
  assign new_n2877_ = ~new_n2876_;
  assign new_n2878_ = new_n2877_ & new_n2875_;
  assign new_n2879_ = new_n2878_ & new_n2873_;
  assign new_n2880_ = ~new_n2879_;
  assign new_n2881_ = new_n2880_ & new_n369_;
  assign new_n2882_ = ~new_n2881_;
  assign new_n2883_ = new_n2882_ & new_n2868_;
  assign new_n2884_ = new_n2883_ & new_n2854_;
  assign new_n2885_ = ~new_n2884_;
  assign new_n2886_ = new_n2885_ & shift6;
  assign new_n2887_ = ~new_n2886_;
  assign new_n2888_ = new_n2887_ & new_n2825_;
  assign ores5 = ~new_n2888_;
  assign new_n2890_ = new_n1859_ & new_n267_;
  assign new_n2891_ = ~new_n2890_;
  assign new_n2892_ = new_n1810_ & new_n293_;
  assign new_n2893_ = ~new_n2892_;
  assign new_n2894_ = new_n2893_ & new_n2891_;
  assign new_n2895_ = new_n1832_ & new_n318_;
  assign new_n2896_ = ~new_n2895_;
  assign new_n2897_ = new_n1817_ & new_n342_;
  assign new_n2898_ = ~new_n2897_;
  assign new_n2899_ = new_n2898_ & new_n2896_;
  assign new_n2900_ = new_n2899_ & new_n2894_;
  assign new_n2901_ = ~new_n2900_;
  assign new_n2902_ = new_n2901_ & new_n369_;
  assign new_n2903_ = ~new_n2902_;
  assign new_n2904_ = new_n1928_ & new_n267_;
  assign new_n2905_ = ~new_n2904_;
  assign new_n2906_ = new_n1844_ & new_n293_;
  assign new_n2907_ = ~new_n2906_;
  assign new_n2908_ = new_n2907_ & new_n2905_;
  assign new_n2909_ = new_n1866_ & new_n318_;
  assign new_n2910_ = ~new_n2909_;
  assign new_n2911_ = new_n1851_ & new_n342_;
  assign new_n2912_ = ~new_n2911_;
  assign new_n2913_ = new_n2912_ & new_n2910_;
  assign new_n2914_ = new_n2913_ & new_n2908_;
  assign new_n2915_ = ~new_n2914_;
  assign new_n2916_ = new_n2915_ & new_n469_;
  assign new_n2917_ = ~new_n2916_;
  assign new_n2918_ = new_n2917_ & new_n2903_;
  assign new_n2919_ = new_n2001_ & new_n267_;
  assign new_n2920_ = ~new_n2919_;
  assign new_n2921_ = new_n1879_ & new_n293_;
  assign new_n2922_ = ~new_n2921_;
  assign new_n2923_ = new_n2922_ & new_n2920_;
  assign new_n2924_ = new_n1901_ & new_n318_;
  assign new_n2925_ = ~new_n2924_;
  assign new_n2926_ = new_n1886_ & new_n342_;
  assign new_n2927_ = ~new_n2926_;
  assign new_n2928_ = new_n2927_ & new_n2925_;
  assign new_n2929_ = new_n2928_ & new_n2923_;
  assign new_n2930_ = ~new_n2929_;
  assign new_n2931_ = new_n2930_ & new_n570_;
  assign new_n2932_ = ~new_n2931_;
  assign new_n2933_ = new_n1894_ & new_n267_;
  assign new_n2934_ = ~new_n2933_;
  assign new_n2935_ = new_n1913_ & new_n293_;
  assign new_n2936_ = ~new_n2935_;
  assign new_n2937_ = new_n2936_ & new_n2934_;
  assign new_n2938_ = new_n1935_ & new_n318_;
  assign new_n2939_ = ~new_n2938_;
  assign new_n2940_ = new_n1920_ & new_n342_;
  assign new_n2941_ = ~new_n2940_;
  assign new_n2942_ = new_n2941_ & new_n2939_;
  assign new_n2943_ = new_n2942_ & new_n2937_;
  assign new_n2944_ = ~new_n2943_;
  assign new_n2945_ = new_n2944_ & new_n669_;
  assign new_n2946_ = ~new_n2945_;
  assign new_n2947_ = new_n2946_ & new_n2932_;
  assign new_n2948_ = new_n2947_ & new_n2918_;
  assign new_n2949_ = ~new_n2948_;
  assign new_n2950_ = new_n2949_ & new_n264_;
  assign new_n2951_ = ~new_n2950_;
  assign new_n2952_ = new_n1967_ & new_n267_;
  assign new_n2953_ = ~new_n2952_;
  assign new_n2954_ = new_n2021_ & new_n293_;
  assign new_n2955_ = ~new_n2954_;
  assign new_n2956_ = new_n2955_ & new_n2953_;
  assign new_n2957_ = new_n2051_ & new_n318_;
  assign new_n2958_ = ~new_n2957_;
  assign new_n2959_ = new_n2028_ & new_n342_;
  assign new_n2960_ = ~new_n2959_;
  assign new_n2961_ = new_n2960_ & new_n2958_;
  assign new_n2962_ = new_n2961_ & new_n2956_;
  assign new_n2963_ = ~new_n2962_;
  assign new_n2964_ = new_n2963_ & new_n669_;
  assign new_n2965_ = ~new_n2964_;
  assign new_n2966_ = new_n1825_ & new_n267_;
  assign new_n2967_ = ~new_n2966_;
  assign new_n2968_ = new_n1952_ & new_n293_;
  assign new_n2969_ = ~new_n2968_;
  assign new_n2970_ = new_n2969_ & new_n2967_;
  assign new_n2971_ = new_n1974_ & new_n318_;
  assign new_n2972_ = ~new_n2971_;
  assign new_n2973_ = new_n1959_ & new_n342_;
  assign new_n2974_ = ~new_n2973_;
  assign new_n2975_ = new_n2974_ & new_n2972_;
  assign new_n2976_ = new_n2975_ & new_n2970_;
  assign new_n2977_ = ~new_n2976_;
  assign new_n2978_ = new_n2977_ & new_n570_;
  assign new_n2979_ = ~new_n2978_;
  assign new_n2980_ = new_n2979_ & new_n2965_;
  assign new_n2981_ = new_n2040_ & new_n267_;
  assign new_n2982_ = ~new_n2981_;
  assign new_n2983_ = new_n2063_ & new_n293_;
  assign new_n2984_ = ~new_n2983_;
  assign new_n2985_ = new_n2984_ & new_n2982_;
  assign new_n2986_ = new_n2085_ & new_n318_;
  assign new_n2987_ = ~new_n2986_;
  assign new_n2988_ = new_n2070_ & new_n342_;
  assign new_n2989_ = ~new_n2988_;
  assign new_n2990_ = new_n2989_ & new_n2987_;
  assign new_n2991_ = new_n2990_ & new_n2985_;
  assign new_n2992_ = ~new_n2991_;
  assign new_n2993_ = new_n2992_ & new_n469_;
  assign new_n2994_ = ~new_n2993_;
  assign new_n2995_ = new_n2078_ & new_n267_;
  assign new_n2996_ = ~new_n2995_;
  assign new_n2997_ = new_n1986_ & new_n293_;
  assign new_n2998_ = ~new_n2997_;
  assign new_n2999_ = new_n2998_ & new_n2996_;
  assign new_n3000_ = new_n2008_ & new_n318_;
  assign new_n3001_ = ~new_n3000_;
  assign new_n3002_ = new_n1993_ & new_n342_;
  assign new_n3003_ = ~new_n3002_;
  assign new_n3004_ = new_n3003_ & new_n3001_;
  assign new_n3005_ = new_n3004_ & new_n2999_;
  assign new_n3006_ = ~new_n3005_;
  assign new_n3007_ = new_n3006_ & new_n369_;
  assign new_n3008_ = ~new_n3007_;
  assign new_n3009_ = new_n3008_ & new_n2994_;
  assign new_n3010_ = new_n3009_ & new_n2980_;
  assign new_n3011_ = ~new_n3010_;
  assign new_n3012_ = new_n3011_ & shift6;
  assign new_n3013_ = ~new_n3012_;
  assign new_n3014_ = new_n3013_ & new_n2951_;
  assign ores6 = ~new_n3014_;
  assign new_n3016_ = new_n2209_ & new_n267_;
  assign new_n3017_ = ~new_n3016_;
  assign new_n3018_ = new_n2311_ & new_n293_;
  assign new_n3019_ = ~new_n3018_;
  assign new_n3020_ = new_n3019_ & new_n3017_;
  assign new_n3021_ = new_n2357_ & new_n318_;
  assign new_n3022_ = ~new_n3021_;
  assign new_n3023_ = new_n2326_ & new_n342_;
  assign new_n3024_ = ~new_n3023_;
  assign new_n3025_ = new_n3024_ & new_n3022_;
  assign new_n3026_ = new_n3025_ & new_n3020_;
  assign new_n3027_ = ~new_n3026_;
  assign new_n3028_ = new_n3027_ & new_n369_;
  assign new_n3029_ = ~new_n3028_;
  assign new_n3030_ = new_n2143_ & new_n267_;
  assign new_n3031_ = ~new_n3030_;
  assign new_n3032_ = new_n2178_ & new_n293_;
  assign new_n3033_ = ~new_n3032_;
  assign new_n3034_ = new_n3033_ & new_n3031_;
  assign new_n3035_ = new_n2224_ & new_n318_;
  assign new_n3036_ = ~new_n3035_;
  assign new_n3037_ = new_n2193_ & new_n342_;
  assign new_n3038_ = ~new_n3037_;
  assign new_n3039_ = new_n3038_ & new_n3036_;
  assign new_n3040_ = new_n3039_ & new_n3034_;
  assign new_n3041_ = ~new_n3040_;
  assign new_n3042_ = new_n3041_ & new_n469_;
  assign new_n3043_ = ~new_n3042_;
  assign new_n3044_ = new_n3043_ & new_n3029_;
  assign new_n3045_ = new_n2542_ & new_n267_;
  assign new_n3046_ = ~new_n3045_;
  assign new_n3047_ = new_n2245_ & new_n293_;
  assign new_n3048_ = ~new_n3047_;
  assign new_n3049_ = new_n3048_ & new_n3046_;
  assign new_n3050_ = new_n2291_ & new_n318_;
  assign new_n3051_ = ~new_n3050_;
  assign new_n3052_ = new_n2260_ & new_n342_;
  assign new_n3053_ = ~new_n3052_;
  assign new_n3054_ = new_n3053_ & new_n3051_;
  assign new_n3055_ = new_n3054_ & new_n3049_;
  assign new_n3056_ = ~new_n3055_;
  assign new_n3057_ = new_n3056_ & new_n570_;
  assign new_n3058_ = ~new_n3057_;
  assign new_n3059_ = new_n2276_ & new_n267_;
  assign new_n3060_ = ~new_n3059_;
  assign new_n3061_ = new_n2112_ & new_n293_;
  assign new_n3062_ = ~new_n3061_;
  assign new_n3063_ = new_n3062_ & new_n3060_;
  assign new_n3064_ = new_n2158_ & new_n318_;
  assign new_n3065_ = ~new_n3064_;
  assign new_n3066_ = new_n2127_ & new_n342_;
  assign new_n3067_ = ~new_n3066_;
  assign new_n3068_ = new_n3067_ & new_n3065_;
  assign new_n3069_ = new_n3068_ & new_n3063_;
  assign new_n3070_ = ~new_n3069_;
  assign new_n3071_ = new_n3070_ & new_n669_;
  assign new_n3072_ = ~new_n3071_;
  assign new_n3073_ = new_n3072_ & new_n3058_;
  assign new_n3074_ = new_n3073_ & new_n3044_;
  assign new_n3075_ = ~new_n3074_;
  assign new_n3076_ = new_n3075_ & new_n264_;
  assign new_n3077_ = ~new_n3076_;
  assign new_n3078_ = new_n2448_ & new_n293_;
  assign new_n3079_ = ~new_n3078_;
  assign new_n3080_ = new_n2459_ & new_n342_;
  assign new_n3081_ = ~new_n3080_;
  assign new_n3082_ = new_n3081_ & new_n3079_;
  assign new_n3083_ = new_n2490_ & new_n318_;
  assign new_n3084_ = ~new_n3083_;
  assign new_n3085_ = new_n2413_ & new_n267_;
  assign new_n3086_ = ~new_n3085_;
  assign new_n3087_ = new_n3086_ & new_n3084_;
  assign new_n3088_ = new_n3087_ & new_n3082_;
  assign new_n3089_ = ~new_n3088_;
  assign new_n3090_ = new_n3089_ & new_n669_;
  assign new_n3091_ = ~new_n3090_;
  assign new_n3092_ = new_n2342_ & new_n267_;
  assign new_n3093_ = ~new_n3092_;
  assign new_n3094_ = new_n2382_ & new_n293_;
  assign new_n3095_ = ~new_n3094_;
  assign new_n3096_ = new_n3095_ & new_n3093_;
  assign new_n3097_ = new_n2428_ & new_n318_;
  assign new_n3098_ = ~new_n3097_;
  assign new_n3099_ = new_n2397_ & new_n342_;
  assign new_n3100_ = ~new_n3099_;
  assign new_n3101_ = new_n3100_ & new_n3098_;
  assign new_n3102_ = new_n3101_ & new_n3096_;
  assign new_n3103_ = ~new_n3102_;
  assign new_n3104_ = new_n3103_ & new_n570_;
  assign new_n3105_ = ~new_n3104_;
  assign new_n3106_ = new_n3105_ & new_n3091_;
  assign new_n3107_ = new_n2475_ & new_n267_;
  assign new_n3108_ = ~new_n3107_;
  assign new_n3109_ = new_n2577_ & new_n293_;
  assign new_n3110_ = ~new_n3109_;
  assign new_n3111_ = new_n3110_ & new_n3108_;
  assign new_n3112_ = new_n2623_ & new_n318_;
  assign new_n3113_ = ~new_n3112_;
  assign new_n3114_ = new_n2592_ & new_n342_;
  assign new_n3115_ = ~new_n3114_;
  assign new_n3116_ = new_n3115_ & new_n3113_;
  assign new_n3117_ = new_n3116_ & new_n3111_;
  assign new_n3118_ = ~new_n3117_;
  assign new_n3119_ = new_n3118_ & new_n469_;
  assign new_n3120_ = ~new_n3119_;
  assign new_n3121_ = new_n2608_ & new_n267_;
  assign new_n3122_ = ~new_n3121_;
  assign new_n3123_ = new_n2511_ & new_n293_;
  assign new_n3124_ = ~new_n3123_;
  assign new_n3125_ = new_n3124_ & new_n3122_;
  assign new_n3126_ = new_n2557_ & new_n318_;
  assign new_n3127_ = ~new_n3126_;
  assign new_n3128_ = new_n2526_ & new_n342_;
  assign new_n3129_ = ~new_n3128_;
  assign new_n3130_ = new_n3129_ & new_n3127_;
  assign new_n3131_ = new_n3130_ & new_n3125_;
  assign new_n3132_ = ~new_n3131_;
  assign new_n3133_ = new_n3132_ & new_n369_;
  assign new_n3134_ = ~new_n3133_;
  assign new_n3135_ = new_n3134_ & new_n3120_;
  assign new_n3136_ = new_n3135_ & new_n3106_;
  assign new_n3137_ = ~new_n3136_;
  assign new_n3138_ = new_n3137_ & shift6;
  assign new_n3139_ = ~new_n3138_;
  assign new_n3140_ = new_n3139_ & new_n3077_;
  assign ores7 = ~new_n3140_;
  assign new_n3142_ = new_n462_ & new_n267_;
  assign new_n3143_ = ~new_n3142_;
  assign new_n3144_ = new_n439_ & new_n293_;
  assign new_n3145_ = ~new_n3144_;
  assign new_n3146_ = new_n3145_ & new_n3143_;
  assign new_n3147_ = new_n318_ & new_n314_;
  assign new_n3148_ = ~new_n3147_;
  assign new_n3149_ = new_n342_ & new_n290_;
  assign new_n3150_ = ~new_n3149_;
  assign new_n3151_ = new_n3150_ & new_n3148_;
  assign new_n3152_ = new_n3151_ & new_n3146_;
  assign new_n3153_ = ~new_n3152_;
  assign new_n3154_ = new_n3153_ & new_n369_;
  assign new_n3155_ = ~new_n3154_;
  assign new_n3156_ = new_n663_ & new_n267_;
  assign new_n3157_ = ~new_n3156_;
  assign new_n3158_ = new_n640_ & new_n293_;
  assign new_n3159_ = ~new_n3158_;
  assign new_n3160_ = new_n3159_ & new_n3157_;
  assign new_n3161_ = new_n415_ & new_n318_;
  assign new_n3162_ = ~new_n3161_;
  assign new_n3163_ = new_n392_ & new_n342_;
  assign new_n3164_ = ~new_n3163_;
  assign new_n3165_ = new_n3164_ & new_n3162_;
  assign new_n3166_ = new_n3165_ & new_n3160_;
  assign new_n3167_ = ~new_n3166_;
  assign new_n3168_ = new_n3167_ & new_n469_;
  assign new_n3169_ = ~new_n3168_;
  assign new_n3170_ = new_n3169_ & new_n3155_;
  assign new_n3171_ = new_n767_ & new_n267_;
  assign new_n3172_ = ~new_n3171_;
  assign new_n3173_ = new_n744_ & new_n293_;
  assign new_n3174_ = ~new_n3173_;
  assign new_n3175_ = new_n3174_ & new_n3172_;
  assign new_n3176_ = new_n516_ & new_n318_;
  assign new_n3177_ = ~new_n3176_;
  assign new_n3178_ = new_n493_ & new_n342_;
  assign new_n3179_ = ~new_n3178_;
  assign new_n3180_ = new_n3179_ & new_n3177_;
  assign new_n3181_ = new_n3180_ & new_n3175_;
  assign new_n3182_ = ~new_n3181_;
  assign new_n3183_ = new_n3182_ & new_n570_;
  assign new_n3184_ = ~new_n3183_;
  assign new_n3185_ = new_n563_ & new_n267_;
  assign new_n3186_ = ~new_n3185_;
  assign new_n3187_ = new_n540_ & new_n293_;
  assign new_n3188_ = ~new_n3187_;
  assign new_n3189_ = new_n3188_ & new_n3186_;
  assign new_n3190_ = new_n616_ & new_n318_;
  assign new_n3191_ = ~new_n3190_;
  assign new_n3192_ = new_n593_ & new_n342_;
  assign new_n3193_ = ~new_n3192_;
  assign new_n3194_ = new_n3193_ & new_n3191_;
  assign new_n3195_ = new_n3194_ & new_n3189_;
  assign new_n3196_ = ~new_n3195_;
  assign new_n3197_ = new_n3196_ & new_n669_;
  assign new_n3198_ = ~new_n3197_;
  assign new_n3199_ = new_n3198_ & new_n3184_;
  assign new_n3200_ = new_n3199_ & new_n3170_;
  assign new_n3201_ = ~new_n3200_;
  assign new_n3202_ = new_n3201_ & new_n264_;
  assign new_n3203_ = ~new_n3202_;
  assign new_n3204_ = new_n964_ & new_n267_;
  assign new_n3205_ = ~new_n3204_;
  assign new_n3206_ = new_n941_ & new_n293_;
  assign new_n3207_ = ~new_n3206_;
  assign new_n3208_ = new_n3207_ & new_n3205_;
  assign new_n3209_ = new_n1015_ & new_n318_;
  assign new_n3210_ = ~new_n3209_;
  assign new_n3211_ = new_n992_ & new_n342_;
  assign new_n3212_ = ~new_n3211_;
  assign new_n3213_ = new_n3212_ & new_n3210_;
  assign new_n3214_ = new_n3213_ & new_n3208_;
  assign new_n3215_ = ~new_n3214_;
  assign new_n3216_ = new_n3215_ & new_n669_;
  assign new_n3217_ = ~new_n3216_;
  assign new_n3218_ = new_n363_ & new_n267_;
  assign new_n3219_ = ~new_n3218_;
  assign new_n3220_ = new_n339_ & new_n293_;
  assign new_n3221_ = ~new_n3220_;
  assign new_n3222_ = new_n3221_ & new_n3219_;
  assign new_n3223_ = new_n917_ & new_n318_;
  assign new_n3224_ = ~new_n3223_;
  assign new_n3225_ = new_n894_ & new_n342_;
  assign new_n3226_ = ~new_n3225_;
  assign new_n3227_ = new_n3226_ & new_n3224_;
  assign new_n3228_ = new_n3227_ & new_n3222_;
  assign new_n3229_ = ~new_n3228_;
  assign new_n3230_ = new_n3229_ & new_n570_;
  assign new_n3231_ = ~new_n3230_;
  assign new_n3232_ = new_n3231_ & new_n3217_;
  assign new_n3233_ = new_n1060_ & new_n267_;
  assign new_n3234_ = ~new_n3233_;
  assign new_n3235_ = new_n1039_ & new_n293_;
  assign new_n3236_ = ~new_n3235_;
  assign new_n3237_ = new_n3236_ & new_n3234_;
  assign new_n3238_ = new_n818_ & new_n318_;
  assign new_n3239_ = ~new_n3238_;
  assign new_n3240_ = new_n795_ & new_n342_;
  assign new_n3241_ = ~new_n3240_;
  assign new_n3242_ = new_n3241_ & new_n3239_;
  assign new_n3243_ = new_n3242_ & new_n3237_;
  assign new_n3244_ = ~new_n3243_;
  assign new_n3245_ = new_n3244_ & new_n469_;
  assign new_n3246_ = ~new_n3245_;
  assign new_n3247_ = new_n865_ & new_n267_;
  assign new_n3248_ = ~new_n3247_;
  assign new_n3249_ = new_n842_ & new_n293_;
  assign new_n3250_ = ~new_n3249_;
  assign new_n3251_ = new_n3250_ & new_n3248_;
  assign new_n3252_ = new_n720_ & new_n318_;
  assign new_n3253_ = ~new_n3252_;
  assign new_n3254_ = new_n697_ & new_n342_;
  assign new_n3255_ = ~new_n3254_;
  assign new_n3256_ = new_n3255_ & new_n3253_;
  assign new_n3257_ = new_n3256_ & new_n3251_;
  assign new_n3258_ = ~new_n3257_;
  assign new_n3259_ = new_n3258_ & new_n369_;
  assign new_n3260_ = ~new_n3259_;
  assign new_n3261_ = new_n3260_ & new_n3246_;
  assign new_n3262_ = new_n3261_ & new_n3232_;
  assign new_n3263_ = ~new_n3262_;
  assign new_n3264_ = new_n3263_ & shift6;
  assign new_n3265_ = ~new_n3264_;
  assign new_n3266_ = new_n3265_ & new_n3203_;
  assign ores8 = ~new_n3266_;
  assign new_n3268_ = new_n1247_ & new_n267_;
  assign new_n3269_ = ~new_n3268_;
  assign new_n3270_ = new_n1226_ & new_n293_;
  assign new_n3271_ = ~new_n3270_;
  assign new_n3272_ = new_n3271_ & new_n3269_;
  assign new_n3273_ = new_n1114_ & new_n318_;
  assign new_n3274_ = ~new_n3273_;
  assign new_n3275_ = new_n1093_ & new_n342_;
  assign new_n3276_ = ~new_n3275_;
  assign new_n3277_ = new_n3276_ & new_n3274_;
  assign new_n3278_ = new_n3277_ & new_n3272_;
  assign new_n3279_ = ~new_n3278_;
  assign new_n3280_ = new_n3279_ & new_n369_;
  assign new_n3281_ = ~new_n3280_;
  assign new_n3282_ = new_n1428_ & new_n267_;
  assign new_n3283_ = ~new_n3282_;
  assign new_n3284_ = new_n1407_ & new_n293_;
  assign new_n3285_ = ~new_n3284_;
  assign new_n3286_ = new_n3285_ & new_n3283_;
  assign new_n3287_ = new_n1204_ & new_n318_;
  assign new_n3288_ = ~new_n3287_;
  assign new_n3289_ = new_n1183_ & new_n342_;
  assign new_n3290_ = ~new_n3289_;
  assign new_n3291_ = new_n3290_ & new_n3288_;
  assign new_n3292_ = new_n3291_ & new_n3286_;
  assign new_n3293_ = ~new_n3292_;
  assign new_n3294_ = new_n3293_ & new_n469_;
  assign new_n3295_ = ~new_n3294_;
  assign new_n3296_ = new_n3295_ & new_n3281_;
  assign new_n3297_ = new_n1613_ & new_n267_;
  assign new_n3298_ = ~new_n3297_;
  assign new_n3299_ = new_n1592_ & new_n293_;
  assign new_n3300_ = ~new_n3299_;
  assign new_n3301_ = new_n3300_ & new_n3298_;
  assign new_n3302_ = new_n1295_ & new_n318_;
  assign new_n3303_ = ~new_n3302_;
  assign new_n3304_ = new_n1274_ & new_n342_;
  assign new_n3305_ = ~new_n3304_;
  assign new_n3306_ = new_n3305_ & new_n3303_;
  assign new_n3307_ = new_n3306_ & new_n3301_;
  assign new_n3308_ = ~new_n3307_;
  assign new_n3309_ = new_n3308_ & new_n570_;
  assign new_n3310_ = ~new_n3309_;
  assign new_n3311_ = new_n1338_ & new_n267_;
  assign new_n3312_ = ~new_n3311_;
  assign new_n3313_ = new_n1317_ & new_n293_;
  assign new_n3314_ = ~new_n3313_;
  assign new_n3315_ = new_n3314_ & new_n3312_;
  assign new_n3316_ = new_n1385_ & new_n318_;
  assign new_n3317_ = ~new_n3316_;
  assign new_n3318_ = new_n1364_ & new_n342_;
  assign new_n3319_ = ~new_n3318_;
  assign new_n3320_ = new_n3319_ & new_n3317_;
  assign new_n3321_ = new_n3320_ & new_n3315_;
  assign new_n3322_ = ~new_n3321_;
  assign new_n3323_ = new_n3322_ & new_n669_;
  assign new_n3324_ = ~new_n3323_;
  assign new_n3325_ = new_n3324_ & new_n3310_;
  assign new_n3326_ = new_n3325_ & new_n3296_;
  assign new_n3327_ = ~new_n3326_;
  assign new_n3328_ = new_n3327_ & new_n264_;
  assign new_n3329_ = ~new_n3328_;
  assign new_n3330_ = new_n1523_ & new_n267_;
  assign new_n3331_ = ~new_n3330_;
  assign new_n3332_ = new_n1502_ & new_n293_;
  assign new_n3333_ = ~new_n3332_;
  assign new_n3334_ = new_n3333_ & new_n3331_;
  assign new_n3335_ = new_n1659_ & new_n318_;
  assign new_n3336_ = ~new_n3335_;
  assign new_n3337_ = new_n1640_ & new_n342_;
  assign new_n3338_ = ~new_n3337_;
  assign new_n3339_ = new_n3338_ & new_n3336_;
  assign new_n3340_ = new_n3339_ & new_n3334_;
  assign new_n3341_ = ~new_n3340_;
  assign new_n3342_ = new_n3341_ & new_n669_;
  assign new_n3343_ = ~new_n3342_;
  assign new_n3344_ = new_n1157_ & new_n267_;
  assign new_n3345_ = ~new_n3344_;
  assign new_n3346_ = new_n1136_ & new_n293_;
  assign new_n3347_ = ~new_n3346_;
  assign new_n3348_ = new_n3347_ & new_n3345_;
  assign new_n3349_ = new_n1480_ & new_n318_;
  assign new_n3350_ = ~new_n3349_;
  assign new_n3351_ = new_n1459_ & new_n342_;
  assign new_n3352_ = ~new_n3351_;
  assign new_n3353_ = new_n3352_ & new_n3350_;
  assign new_n3354_ = new_n3353_ & new_n3348_;
  assign new_n3355_ = ~new_n3354_;
  assign new_n3356_ = new_n3355_ & new_n570_;
  assign new_n3357_ = ~new_n3356_;
  assign new_n3358_ = new_n3357_ & new_n3343_;
  assign new_n3359_ = new_n1701_ & new_n267_;
  assign new_n3360_ = ~new_n3359_;
  assign new_n3361_ = new_n1681_ & new_n293_;
  assign new_n3362_ = ~new_n3361_;
  assign new_n3363_ = new_n3362_ & new_n3360_;
  assign new_n3364_ = new_n1748_ & new_n318_;
  assign new_n3365_ = ~new_n3364_;
  assign new_n3366_ = new_n1727_ & new_n342_;
  assign new_n3367_ = ~new_n3366_;
  assign new_n3368_ = new_n3367_ & new_n3365_;
  assign new_n3369_ = new_n3368_ & new_n3363_;
  assign new_n3370_ = ~new_n3369_;
  assign new_n3371_ = new_n3370_ & new_n469_;
  assign new_n3372_ = ~new_n3371_;
  assign new_n3373_ = new_n1791_ & new_n267_;
  assign new_n3374_ = ~new_n3373_;
  assign new_n3375_ = new_n1770_ & new_n293_;
  assign new_n3376_ = ~new_n3375_;
  assign new_n3377_ = new_n3376_ & new_n3374_;
  assign new_n3378_ = new_n1570_ & new_n318_;
  assign new_n3379_ = ~new_n3378_;
  assign new_n3380_ = new_n1549_ & new_n342_;
  assign new_n3381_ = ~new_n3380_;
  assign new_n3382_ = new_n3381_ & new_n3379_;
  assign new_n3383_ = new_n3382_ & new_n3377_;
  assign new_n3384_ = ~new_n3383_;
  assign new_n3385_ = new_n3384_ & new_n369_;
  assign new_n3386_ = ~new_n3385_;
  assign new_n3387_ = new_n3386_ & new_n3372_;
  assign new_n3388_ = new_n3387_ & new_n3358_;
  assign new_n3389_ = ~new_n3388_;
  assign new_n3390_ = new_n3389_ & shift6;
  assign new_n3391_ = ~new_n3390_;
  assign new_n3392_ = new_n3391_ & new_n3329_;
  assign ores9 = ~new_n3392_;
  assign new_n3394_ = new_n1866_ & new_n267_;
  assign new_n3395_ = ~new_n3394_;
  assign new_n3396_ = new_n1859_ & new_n293_;
  assign new_n3397_ = ~new_n3396_;
  assign new_n3398_ = new_n3397_ & new_n3395_;
  assign new_n3399_ = new_n1817_ & new_n318_;
  assign new_n3400_ = ~new_n3399_;
  assign new_n3401_ = new_n1810_ & new_n342_;
  assign new_n3402_ = ~new_n3401_;
  assign new_n3403_ = new_n3402_ & new_n3400_;
  assign new_n3404_ = new_n3403_ & new_n3398_;
  assign new_n3405_ = ~new_n3404_;
  assign new_n3406_ = new_n3405_ & new_n369_;
  assign new_n3407_ = ~new_n3406_;
  assign new_n3408_ = new_n1935_ & new_n267_;
  assign new_n3409_ = ~new_n3408_;
  assign new_n3410_ = new_n1928_ & new_n293_;
  assign new_n3411_ = ~new_n3410_;
  assign new_n3412_ = new_n3411_ & new_n3409_;
  assign new_n3413_ = new_n1851_ & new_n318_;
  assign new_n3414_ = ~new_n3413_;
  assign new_n3415_ = new_n1844_ & new_n342_;
  assign new_n3416_ = ~new_n3415_;
  assign new_n3417_ = new_n3416_ & new_n3414_;
  assign new_n3418_ = new_n3417_ & new_n3412_;
  assign new_n3419_ = ~new_n3418_;
  assign new_n3420_ = new_n3419_ & new_n469_;
  assign new_n3421_ = ~new_n3420_;
  assign new_n3422_ = new_n3421_ & new_n3407_;
  assign new_n3423_ = new_n2008_ & new_n267_;
  assign new_n3424_ = ~new_n3423_;
  assign new_n3425_ = new_n2001_ & new_n293_;
  assign new_n3426_ = ~new_n3425_;
  assign new_n3427_ = new_n3426_ & new_n3424_;
  assign new_n3428_ = new_n1886_ & new_n318_;
  assign new_n3429_ = ~new_n3428_;
  assign new_n3430_ = new_n1879_ & new_n342_;
  assign new_n3431_ = ~new_n3430_;
  assign new_n3432_ = new_n3431_ & new_n3429_;
  assign new_n3433_ = new_n3432_ & new_n3427_;
  assign new_n3434_ = ~new_n3433_;
  assign new_n3435_ = new_n3434_ & new_n570_;
  assign new_n3436_ = ~new_n3435_;
  assign new_n3437_ = new_n1901_ & new_n267_;
  assign new_n3438_ = ~new_n3437_;
  assign new_n3439_ = new_n1894_ & new_n293_;
  assign new_n3440_ = ~new_n3439_;
  assign new_n3441_ = new_n3440_ & new_n3438_;
  assign new_n3442_ = new_n1920_ & new_n318_;
  assign new_n3443_ = ~new_n3442_;
  assign new_n3444_ = new_n1913_ & new_n342_;
  assign new_n3445_ = ~new_n3444_;
  assign new_n3446_ = new_n3445_ & new_n3443_;
  assign new_n3447_ = new_n3446_ & new_n3441_;
  assign new_n3448_ = ~new_n3447_;
  assign new_n3449_ = new_n3448_ & new_n669_;
  assign new_n3450_ = ~new_n3449_;
  assign new_n3451_ = new_n3450_ & new_n3436_;
  assign new_n3452_ = new_n3451_ & new_n3422_;
  assign new_n3453_ = ~new_n3452_;
  assign new_n3454_ = new_n3453_ & new_n264_;
  assign new_n3455_ = ~new_n3454_;
  assign new_n3456_ = new_n1974_ & new_n267_;
  assign new_n3457_ = ~new_n3456_;
  assign new_n3458_ = new_n1967_ & new_n293_;
  assign new_n3459_ = ~new_n3458_;
  assign new_n3460_ = new_n3459_ & new_n3457_;
  assign new_n3461_ = new_n2028_ & new_n318_;
  assign new_n3462_ = ~new_n3461_;
  assign new_n3463_ = new_n2021_ & new_n342_;
  assign new_n3464_ = ~new_n3463_;
  assign new_n3465_ = new_n3464_ & new_n3462_;
  assign new_n3466_ = new_n3465_ & new_n3460_;
  assign new_n3467_ = ~new_n3466_;
  assign new_n3468_ = new_n3467_ & new_n669_;
  assign new_n3469_ = ~new_n3468_;
  assign new_n3470_ = new_n1832_ & new_n267_;
  assign new_n3471_ = ~new_n3470_;
  assign new_n3472_ = new_n1825_ & new_n293_;
  assign new_n3473_ = ~new_n3472_;
  assign new_n3474_ = new_n3473_ & new_n3471_;
  assign new_n3475_ = new_n1959_ & new_n318_;
  assign new_n3476_ = ~new_n3475_;
  assign new_n3477_ = new_n1952_ & new_n342_;
  assign new_n3478_ = ~new_n3477_;
  assign new_n3479_ = new_n3478_ & new_n3476_;
  assign new_n3480_ = new_n3479_ & new_n3474_;
  assign new_n3481_ = ~new_n3480_;
  assign new_n3482_ = new_n3481_ & new_n570_;
  assign new_n3483_ = ~new_n3482_;
  assign new_n3484_ = new_n3483_ & new_n3469_;
  assign new_n3485_ = new_n2051_ & new_n267_;
  assign new_n3486_ = ~new_n3485_;
  assign new_n3487_ = new_n2040_ & new_n293_;
  assign new_n3488_ = ~new_n3487_;
  assign new_n3489_ = new_n3488_ & new_n3486_;
  assign new_n3490_ = new_n2070_ & new_n318_;
  assign new_n3491_ = ~new_n3490_;
  assign new_n3492_ = new_n2063_ & new_n342_;
  assign new_n3493_ = ~new_n3492_;
  assign new_n3494_ = new_n3493_ & new_n3491_;
  assign new_n3495_ = new_n3494_ & new_n3489_;
  assign new_n3496_ = ~new_n3495_;
  assign new_n3497_ = new_n3496_ & new_n469_;
  assign new_n3498_ = ~new_n3497_;
  assign new_n3499_ = new_n2085_ & new_n267_;
  assign new_n3500_ = ~new_n3499_;
  assign new_n3501_ = new_n2078_ & new_n293_;
  assign new_n3502_ = ~new_n3501_;
  assign new_n3503_ = new_n3502_ & new_n3500_;
  assign new_n3504_ = new_n1993_ & new_n318_;
  assign new_n3505_ = ~new_n3504_;
  assign new_n3506_ = new_n1986_ & new_n342_;
  assign new_n3507_ = ~new_n3506_;
  assign new_n3508_ = new_n3507_ & new_n3505_;
  assign new_n3509_ = new_n3508_ & new_n3503_;
  assign new_n3510_ = ~new_n3509_;
  assign new_n3511_ = new_n3510_ & new_n369_;
  assign new_n3512_ = ~new_n3511_;
  assign new_n3513_ = new_n3512_ & new_n3498_;
  assign new_n3514_ = new_n3513_ & new_n3484_;
  assign new_n3515_ = ~new_n3514_;
  assign new_n3516_ = new_n3515_ & shift6;
  assign new_n3517_ = ~new_n3516_;
  assign new_n3518_ = new_n3517_ & new_n3455_;
  assign ores10 = ~new_n3518_;
  assign new_n3520_ = new_n2224_ & new_n267_;
  assign new_n3521_ = ~new_n3520_;
  assign new_n3522_ = new_n2209_ & new_n293_;
  assign new_n3523_ = ~new_n3522_;
  assign new_n3524_ = new_n3523_ & new_n3521_;
  assign new_n3525_ = new_n2326_ & new_n318_;
  assign new_n3526_ = ~new_n3525_;
  assign new_n3527_ = new_n2311_ & new_n342_;
  assign new_n3528_ = ~new_n3527_;
  assign new_n3529_ = new_n3528_ & new_n3526_;
  assign new_n3530_ = new_n3529_ & new_n3524_;
  assign new_n3531_ = ~new_n3530_;
  assign new_n3532_ = new_n3531_ & new_n369_;
  assign new_n3533_ = ~new_n3532_;
  assign new_n3534_ = new_n2158_ & new_n267_;
  assign new_n3535_ = ~new_n3534_;
  assign new_n3536_ = new_n2143_ & new_n293_;
  assign new_n3537_ = ~new_n3536_;
  assign new_n3538_ = new_n3537_ & new_n3535_;
  assign new_n3539_ = new_n2193_ & new_n318_;
  assign new_n3540_ = ~new_n3539_;
  assign new_n3541_ = new_n2178_ & new_n342_;
  assign new_n3542_ = ~new_n3541_;
  assign new_n3543_ = new_n3542_ & new_n3540_;
  assign new_n3544_ = new_n3543_ & new_n3538_;
  assign new_n3545_ = ~new_n3544_;
  assign new_n3546_ = new_n3545_ & new_n469_;
  assign new_n3547_ = ~new_n3546_;
  assign new_n3548_ = new_n3547_ & new_n3533_;
  assign new_n3549_ = new_n2557_ & new_n267_;
  assign new_n3550_ = ~new_n3549_;
  assign new_n3551_ = new_n2542_ & new_n293_;
  assign new_n3552_ = ~new_n3551_;
  assign new_n3553_ = new_n3552_ & new_n3550_;
  assign new_n3554_ = new_n2260_ & new_n318_;
  assign new_n3555_ = ~new_n3554_;
  assign new_n3556_ = new_n2245_ & new_n342_;
  assign new_n3557_ = ~new_n3556_;
  assign new_n3558_ = new_n3557_ & new_n3555_;
  assign new_n3559_ = new_n3558_ & new_n3553_;
  assign new_n3560_ = ~new_n3559_;
  assign new_n3561_ = new_n3560_ & new_n570_;
  assign new_n3562_ = ~new_n3561_;
  assign new_n3563_ = new_n2291_ & new_n267_;
  assign new_n3564_ = ~new_n3563_;
  assign new_n3565_ = new_n2276_ & new_n293_;
  assign new_n3566_ = ~new_n3565_;
  assign new_n3567_ = new_n3566_ & new_n3564_;
  assign new_n3568_ = new_n2127_ & new_n318_;
  assign new_n3569_ = ~new_n3568_;
  assign new_n3570_ = new_n2112_ & new_n342_;
  assign new_n3571_ = ~new_n3570_;
  assign new_n3572_ = new_n3571_ & new_n3569_;
  assign new_n3573_ = new_n3572_ & new_n3567_;
  assign new_n3574_ = ~new_n3573_;
  assign new_n3575_ = new_n3574_ & new_n669_;
  assign new_n3576_ = ~new_n3575_;
  assign new_n3577_ = new_n3576_ & new_n3562_;
  assign new_n3578_ = new_n3577_ & new_n3548_;
  assign new_n3579_ = ~new_n3578_;
  assign new_n3580_ = new_n3579_ & new_n264_;
  assign new_n3581_ = ~new_n3580_;
  assign new_n3582_ = new_n2428_ & new_n267_;
  assign new_n3583_ = ~new_n3582_;
  assign new_n3584_ = new_n2448_ & new_n342_;
  assign new_n3585_ = ~new_n3584_;
  assign new_n3586_ = new_n3585_ & new_n3583_;
  assign new_n3587_ = new_n2459_ & new_n318_;
  assign new_n3588_ = ~new_n3587_;
  assign new_n3589_ = new_n2413_ & new_n293_;
  assign new_n3590_ = ~new_n3589_;
  assign new_n3591_ = new_n3590_ & new_n3588_;
  assign new_n3592_ = new_n3591_ & new_n3586_;
  assign new_n3593_ = ~new_n3592_;
  assign new_n3594_ = new_n3593_ & new_n669_;
  assign new_n3595_ = ~new_n3594_;
  assign new_n3596_ = new_n2357_ & new_n267_;
  assign new_n3597_ = ~new_n3596_;
  assign new_n3598_ = new_n2342_ & new_n293_;
  assign new_n3599_ = ~new_n3598_;
  assign new_n3600_ = new_n3599_ & new_n3597_;
  assign new_n3601_ = new_n2397_ & new_n318_;
  assign new_n3602_ = ~new_n3601_;
  assign new_n3603_ = new_n2382_ & new_n342_;
  assign new_n3604_ = ~new_n3603_;
  assign new_n3605_ = new_n3604_ & new_n3602_;
  assign new_n3606_ = new_n3605_ & new_n3600_;
  assign new_n3607_ = ~new_n3606_;
  assign new_n3608_ = new_n3607_ & new_n570_;
  assign new_n3609_ = ~new_n3608_;
  assign new_n3610_ = new_n3609_ & new_n3595_;
  assign new_n3611_ = new_n2490_ & new_n267_;
  assign new_n3612_ = ~new_n3611_;
  assign new_n3613_ = new_n2475_ & new_n293_;
  assign new_n3614_ = ~new_n3613_;
  assign new_n3615_ = new_n3614_ & new_n3612_;
  assign new_n3616_ = new_n2592_ & new_n318_;
  assign new_n3617_ = ~new_n3616_;
  assign new_n3618_ = new_n2577_ & new_n342_;
  assign new_n3619_ = ~new_n3618_;
  assign new_n3620_ = new_n3619_ & new_n3617_;
  assign new_n3621_ = new_n3620_ & new_n3615_;
  assign new_n3622_ = ~new_n3621_;
  assign new_n3623_ = new_n3622_ & new_n469_;
  assign new_n3624_ = ~new_n3623_;
  assign new_n3625_ = new_n2623_ & new_n267_;
  assign new_n3626_ = ~new_n3625_;
  assign new_n3627_ = new_n2608_ & new_n293_;
  assign new_n3628_ = ~new_n3627_;
  assign new_n3629_ = new_n3628_ & new_n3626_;
  assign new_n3630_ = new_n2526_ & new_n318_;
  assign new_n3631_ = ~new_n3630_;
  assign new_n3632_ = new_n2511_ & new_n342_;
  assign new_n3633_ = ~new_n3632_;
  assign new_n3634_ = new_n3633_ & new_n3631_;
  assign new_n3635_ = new_n3634_ & new_n3629_;
  assign new_n3636_ = ~new_n3635_;
  assign new_n3637_ = new_n3636_ & new_n369_;
  assign new_n3638_ = ~new_n3637_;
  assign new_n3639_ = new_n3638_ & new_n3624_;
  assign new_n3640_ = new_n3639_ & new_n3610_;
  assign new_n3641_ = ~new_n3640_;
  assign new_n3642_ = new_n3641_ & shift6;
  assign new_n3643_ = ~new_n3642_;
  assign new_n3644_ = new_n3643_ & new_n3581_;
  assign ores11 = ~new_n3644_;
  assign new_n3646_ = new_n415_ & new_n267_;
  assign new_n3647_ = ~new_n3646_;
  assign new_n3648_ = new_n462_ & new_n293_;
  assign new_n3649_ = ~new_n3648_;
  assign new_n3650_ = new_n3649_ & new_n3647_;
  assign new_n3651_ = new_n318_ & new_n290_;
  assign new_n3652_ = ~new_n3651_;
  assign new_n3653_ = new_n439_ & new_n342_;
  assign new_n3654_ = ~new_n3653_;
  assign new_n3655_ = new_n3654_ & new_n3652_;
  assign new_n3656_ = new_n3655_ & new_n3650_;
  assign new_n3657_ = ~new_n3656_;
  assign new_n3658_ = new_n3657_ & new_n369_;
  assign new_n3659_ = ~new_n3658_;
  assign new_n3660_ = new_n616_ & new_n267_;
  assign new_n3661_ = ~new_n3660_;
  assign new_n3662_ = new_n663_ & new_n293_;
  assign new_n3663_ = ~new_n3662_;
  assign new_n3664_ = new_n3663_ & new_n3661_;
  assign new_n3665_ = new_n392_ & new_n318_;
  assign new_n3666_ = ~new_n3665_;
  assign new_n3667_ = new_n640_ & new_n342_;
  assign new_n3668_ = ~new_n3667_;
  assign new_n3669_ = new_n3668_ & new_n3666_;
  assign new_n3670_ = new_n3669_ & new_n3664_;
  assign new_n3671_ = ~new_n3670_;
  assign new_n3672_ = new_n3671_ & new_n469_;
  assign new_n3673_ = ~new_n3672_;
  assign new_n3674_ = new_n3673_ & new_n3659_;
  assign new_n3675_ = new_n720_ & new_n267_;
  assign new_n3676_ = ~new_n3675_;
  assign new_n3677_ = new_n767_ & new_n293_;
  assign new_n3678_ = ~new_n3677_;
  assign new_n3679_ = new_n3678_ & new_n3676_;
  assign new_n3680_ = new_n493_ & new_n318_;
  assign new_n3681_ = ~new_n3680_;
  assign new_n3682_ = new_n744_ & new_n342_;
  assign new_n3683_ = ~new_n3682_;
  assign new_n3684_ = new_n3683_ & new_n3681_;
  assign new_n3685_ = new_n3684_ & new_n3679_;
  assign new_n3686_ = ~new_n3685_;
  assign new_n3687_ = new_n3686_ & new_n570_;
  assign new_n3688_ = ~new_n3687_;
  assign new_n3689_ = new_n516_ & new_n267_;
  assign new_n3690_ = ~new_n3689_;
  assign new_n3691_ = new_n563_ & new_n293_;
  assign new_n3692_ = ~new_n3691_;
  assign new_n3693_ = new_n3692_ & new_n3690_;
  assign new_n3694_ = new_n593_ & new_n318_;
  assign new_n3695_ = ~new_n3694_;
  assign new_n3696_ = new_n540_ & new_n342_;
  assign new_n3697_ = ~new_n3696_;
  assign new_n3698_ = new_n3697_ & new_n3695_;
  assign new_n3699_ = new_n3698_ & new_n3693_;
  assign new_n3700_ = ~new_n3699_;
  assign new_n3701_ = new_n3700_ & new_n669_;
  assign new_n3702_ = ~new_n3701_;
  assign new_n3703_ = new_n3702_ & new_n3688_;
  assign new_n3704_ = new_n3703_ & new_n3674_;
  assign new_n3705_ = ~new_n3704_;
  assign new_n3706_ = new_n3705_ & new_n264_;
  assign new_n3707_ = ~new_n3706_;
  assign new_n3708_ = new_n917_ & new_n267_;
  assign new_n3709_ = ~new_n3708_;
  assign new_n3710_ = new_n964_ & new_n293_;
  assign new_n3711_ = ~new_n3710_;
  assign new_n3712_ = new_n3711_ & new_n3709_;
  assign new_n3713_ = new_n992_ & new_n318_;
  assign new_n3714_ = ~new_n3713_;
  assign new_n3715_ = new_n941_ & new_n342_;
  assign new_n3716_ = ~new_n3715_;
  assign new_n3717_ = new_n3716_ & new_n3714_;
  assign new_n3718_ = new_n3717_ & new_n3712_;
  assign new_n3719_ = ~new_n3718_;
  assign new_n3720_ = new_n3719_ & new_n669_;
  assign new_n3721_ = ~new_n3720_;
  assign new_n3722_ = new_n314_ & new_n267_;
  assign new_n3723_ = ~new_n3722_;
  assign new_n3724_ = new_n363_ & new_n293_;
  assign new_n3725_ = ~new_n3724_;
  assign new_n3726_ = new_n3725_ & new_n3723_;
  assign new_n3727_ = new_n894_ & new_n318_;
  assign new_n3728_ = ~new_n3727_;
  assign new_n3729_ = new_n342_ & new_n339_;
  assign new_n3730_ = ~new_n3729_;
  assign new_n3731_ = new_n3730_ & new_n3728_;
  assign new_n3732_ = new_n3731_ & new_n3726_;
  assign new_n3733_ = ~new_n3732_;
  assign new_n3734_ = new_n3733_ & new_n570_;
  assign new_n3735_ = ~new_n3734_;
  assign new_n3736_ = new_n3735_ & new_n3721_;
  assign new_n3737_ = new_n1015_ & new_n267_;
  assign new_n3738_ = ~new_n3737_;
  assign new_n3739_ = new_n1060_ & new_n293_;
  assign new_n3740_ = ~new_n3739_;
  assign new_n3741_ = new_n3740_ & new_n3738_;
  assign new_n3742_ = new_n795_ & new_n318_;
  assign new_n3743_ = ~new_n3742_;
  assign new_n3744_ = new_n1039_ & new_n342_;
  assign new_n3745_ = ~new_n3744_;
  assign new_n3746_ = new_n3745_ & new_n3743_;
  assign new_n3747_ = new_n3746_ & new_n3741_;
  assign new_n3748_ = ~new_n3747_;
  assign new_n3749_ = new_n3748_ & new_n469_;
  assign new_n3750_ = ~new_n3749_;
  assign new_n3751_ = new_n818_ & new_n267_;
  assign new_n3752_ = ~new_n3751_;
  assign new_n3753_ = new_n865_ & new_n293_;
  assign new_n3754_ = ~new_n3753_;
  assign new_n3755_ = new_n3754_ & new_n3752_;
  assign new_n3756_ = new_n697_ & new_n318_;
  assign new_n3757_ = ~new_n3756_;
  assign new_n3758_ = new_n842_ & new_n342_;
  assign new_n3759_ = ~new_n3758_;
  assign new_n3760_ = new_n3759_ & new_n3757_;
  assign new_n3761_ = new_n3760_ & new_n3755_;
  assign new_n3762_ = ~new_n3761_;
  assign new_n3763_ = new_n3762_ & new_n369_;
  assign new_n3764_ = ~new_n3763_;
  assign new_n3765_ = new_n3764_ & new_n3750_;
  assign new_n3766_ = new_n3765_ & new_n3736_;
  assign new_n3767_ = ~new_n3766_;
  assign new_n3768_ = new_n3767_ & shift6;
  assign new_n3769_ = ~new_n3768_;
  assign new_n3770_ = new_n3769_ & new_n3707_;
  assign ores12 = ~new_n3770_;
  assign new_n3772_ = new_n1204_ & new_n267_;
  assign new_n3773_ = ~new_n3772_;
  assign new_n3774_ = new_n1247_ & new_n293_;
  assign new_n3775_ = ~new_n3774_;
  assign new_n3776_ = new_n3775_ & new_n3773_;
  assign new_n3777_ = new_n1093_ & new_n318_;
  assign new_n3778_ = ~new_n3777_;
  assign new_n3779_ = new_n1226_ & new_n342_;
  assign new_n3780_ = ~new_n3779_;
  assign new_n3781_ = new_n3780_ & new_n3778_;
  assign new_n3782_ = new_n3781_ & new_n3776_;
  assign new_n3783_ = ~new_n3782_;
  assign new_n3784_ = new_n3783_ & new_n369_;
  assign new_n3785_ = ~new_n3784_;
  assign new_n3786_ = new_n1385_ & new_n267_;
  assign new_n3787_ = ~new_n3786_;
  assign new_n3788_ = new_n1428_ & new_n293_;
  assign new_n3789_ = ~new_n3788_;
  assign new_n3790_ = new_n3789_ & new_n3787_;
  assign new_n3791_ = new_n1183_ & new_n318_;
  assign new_n3792_ = ~new_n3791_;
  assign new_n3793_ = new_n1407_ & new_n342_;
  assign new_n3794_ = ~new_n3793_;
  assign new_n3795_ = new_n3794_ & new_n3792_;
  assign new_n3796_ = new_n3795_ & new_n3790_;
  assign new_n3797_ = ~new_n3796_;
  assign new_n3798_ = new_n3797_ & new_n469_;
  assign new_n3799_ = ~new_n3798_;
  assign new_n3800_ = new_n3799_ & new_n3785_;
  assign new_n3801_ = new_n1570_ & new_n267_;
  assign new_n3802_ = ~new_n3801_;
  assign new_n3803_ = new_n1613_ & new_n293_;
  assign new_n3804_ = ~new_n3803_;
  assign new_n3805_ = new_n3804_ & new_n3802_;
  assign new_n3806_ = new_n1274_ & new_n318_;
  assign new_n3807_ = ~new_n3806_;
  assign new_n3808_ = new_n1592_ & new_n342_;
  assign new_n3809_ = ~new_n3808_;
  assign new_n3810_ = new_n3809_ & new_n3807_;
  assign new_n3811_ = new_n3810_ & new_n3805_;
  assign new_n3812_ = ~new_n3811_;
  assign new_n3813_ = new_n3812_ & new_n570_;
  assign new_n3814_ = ~new_n3813_;
  assign new_n3815_ = new_n1295_ & new_n267_;
  assign new_n3816_ = ~new_n3815_;
  assign new_n3817_ = new_n1338_ & new_n293_;
  assign new_n3818_ = ~new_n3817_;
  assign new_n3819_ = new_n3818_ & new_n3816_;
  assign new_n3820_ = new_n1364_ & new_n318_;
  assign new_n3821_ = ~new_n3820_;
  assign new_n3822_ = new_n1317_ & new_n342_;
  assign new_n3823_ = ~new_n3822_;
  assign new_n3824_ = new_n3823_ & new_n3821_;
  assign new_n3825_ = new_n3824_ & new_n3819_;
  assign new_n3826_ = ~new_n3825_;
  assign new_n3827_ = new_n3826_ & new_n669_;
  assign new_n3828_ = ~new_n3827_;
  assign new_n3829_ = new_n3828_ & new_n3814_;
  assign new_n3830_ = new_n3829_ & new_n3800_;
  assign new_n3831_ = ~new_n3830_;
  assign new_n3832_ = new_n3831_ & new_n264_;
  assign new_n3833_ = ~new_n3832_;
  assign new_n3834_ = new_n1480_ & new_n267_;
  assign new_n3835_ = ~new_n3834_;
  assign new_n3836_ = new_n1523_ & new_n293_;
  assign new_n3837_ = ~new_n3836_;
  assign new_n3838_ = new_n3837_ & new_n3835_;
  assign new_n3839_ = new_n1640_ & new_n318_;
  assign new_n3840_ = ~new_n3839_;
  assign new_n3841_ = new_n1502_ & new_n342_;
  assign new_n3842_ = ~new_n3841_;
  assign new_n3843_ = new_n3842_ & new_n3840_;
  assign new_n3844_ = new_n3843_ & new_n3838_;
  assign new_n3845_ = ~new_n3844_;
  assign new_n3846_ = new_n3845_ & new_n669_;
  assign new_n3847_ = ~new_n3846_;
  assign new_n3848_ = new_n1114_ & new_n267_;
  assign new_n3849_ = ~new_n3848_;
  assign new_n3850_ = new_n1157_ & new_n293_;
  assign new_n3851_ = ~new_n3850_;
  assign new_n3852_ = new_n3851_ & new_n3849_;
  assign new_n3853_ = new_n1459_ & new_n318_;
  assign new_n3854_ = ~new_n3853_;
  assign new_n3855_ = new_n1136_ & new_n342_;
  assign new_n3856_ = ~new_n3855_;
  assign new_n3857_ = new_n3856_ & new_n3854_;
  assign new_n3858_ = new_n3857_ & new_n3852_;
  assign new_n3859_ = ~new_n3858_;
  assign new_n3860_ = new_n3859_ & new_n570_;
  assign new_n3861_ = ~new_n3860_;
  assign new_n3862_ = new_n3861_ & new_n3847_;
  assign new_n3863_ = new_n1659_ & new_n267_;
  assign new_n3864_ = ~new_n3863_;
  assign new_n3865_ = new_n1701_ & new_n293_;
  assign new_n3866_ = ~new_n3865_;
  assign new_n3867_ = new_n3866_ & new_n3864_;
  assign new_n3868_ = new_n1727_ & new_n318_;
  assign new_n3869_ = ~new_n3868_;
  assign new_n3870_ = new_n1681_ & new_n342_;
  assign new_n3871_ = ~new_n3870_;
  assign new_n3872_ = new_n3871_ & new_n3869_;
  assign new_n3873_ = new_n3872_ & new_n3867_;
  assign new_n3874_ = ~new_n3873_;
  assign new_n3875_ = new_n3874_ & new_n469_;
  assign new_n3876_ = ~new_n3875_;
  assign new_n3877_ = new_n1748_ & new_n267_;
  assign new_n3878_ = ~new_n3877_;
  assign new_n3879_ = new_n1791_ & new_n293_;
  assign new_n3880_ = ~new_n3879_;
  assign new_n3881_ = new_n3880_ & new_n3878_;
  assign new_n3882_ = new_n1549_ & new_n318_;
  assign new_n3883_ = ~new_n3882_;
  assign new_n3884_ = new_n1770_ & new_n342_;
  assign new_n3885_ = ~new_n3884_;
  assign new_n3886_ = new_n3885_ & new_n3883_;
  assign new_n3887_ = new_n3886_ & new_n3881_;
  assign new_n3888_ = ~new_n3887_;
  assign new_n3889_ = new_n3888_ & new_n369_;
  assign new_n3890_ = ~new_n3889_;
  assign new_n3891_ = new_n3890_ & new_n3876_;
  assign new_n3892_ = new_n3891_ & new_n3862_;
  assign new_n3893_ = ~new_n3892_;
  assign new_n3894_ = new_n3893_ & shift6;
  assign new_n3895_ = ~new_n3894_;
  assign new_n3896_ = new_n3895_ & new_n3833_;
  assign ores13 = ~new_n3896_;
  assign new_n3898_ = new_n1851_ & new_n267_;
  assign new_n3899_ = ~new_n3898_;
  assign new_n3900_ = new_n1866_ & new_n293_;
  assign new_n3901_ = ~new_n3900_;
  assign new_n3902_ = new_n3901_ & new_n3899_;
  assign new_n3903_ = new_n1810_ & new_n318_;
  assign new_n3904_ = ~new_n3903_;
  assign new_n3905_ = new_n1859_ & new_n342_;
  assign new_n3906_ = ~new_n3905_;
  assign new_n3907_ = new_n3906_ & new_n3904_;
  assign new_n3908_ = new_n3907_ & new_n3902_;
  assign new_n3909_ = ~new_n3908_;
  assign new_n3910_ = new_n3909_ & new_n369_;
  assign new_n3911_ = ~new_n3910_;
  assign new_n3912_ = new_n1920_ & new_n267_;
  assign new_n3913_ = ~new_n3912_;
  assign new_n3914_ = new_n1935_ & new_n293_;
  assign new_n3915_ = ~new_n3914_;
  assign new_n3916_ = new_n3915_ & new_n3913_;
  assign new_n3917_ = new_n1844_ & new_n318_;
  assign new_n3918_ = ~new_n3917_;
  assign new_n3919_ = new_n1928_ & new_n342_;
  assign new_n3920_ = ~new_n3919_;
  assign new_n3921_ = new_n3920_ & new_n3918_;
  assign new_n3922_ = new_n3921_ & new_n3916_;
  assign new_n3923_ = ~new_n3922_;
  assign new_n3924_ = new_n3923_ & new_n469_;
  assign new_n3925_ = ~new_n3924_;
  assign new_n3926_ = new_n3925_ & new_n3911_;
  assign new_n3927_ = new_n1993_ & new_n267_;
  assign new_n3928_ = ~new_n3927_;
  assign new_n3929_ = new_n2008_ & new_n293_;
  assign new_n3930_ = ~new_n3929_;
  assign new_n3931_ = new_n3930_ & new_n3928_;
  assign new_n3932_ = new_n1879_ & new_n318_;
  assign new_n3933_ = ~new_n3932_;
  assign new_n3934_ = new_n2001_ & new_n342_;
  assign new_n3935_ = ~new_n3934_;
  assign new_n3936_ = new_n3935_ & new_n3933_;
  assign new_n3937_ = new_n3936_ & new_n3931_;
  assign new_n3938_ = ~new_n3937_;
  assign new_n3939_ = new_n3938_ & new_n570_;
  assign new_n3940_ = ~new_n3939_;
  assign new_n3941_ = new_n1886_ & new_n267_;
  assign new_n3942_ = ~new_n3941_;
  assign new_n3943_ = new_n1901_ & new_n293_;
  assign new_n3944_ = ~new_n3943_;
  assign new_n3945_ = new_n3944_ & new_n3942_;
  assign new_n3946_ = new_n1913_ & new_n318_;
  assign new_n3947_ = ~new_n3946_;
  assign new_n3948_ = new_n1894_ & new_n342_;
  assign new_n3949_ = ~new_n3948_;
  assign new_n3950_ = new_n3949_ & new_n3947_;
  assign new_n3951_ = new_n3950_ & new_n3945_;
  assign new_n3952_ = ~new_n3951_;
  assign new_n3953_ = new_n3952_ & new_n669_;
  assign new_n3954_ = ~new_n3953_;
  assign new_n3955_ = new_n3954_ & new_n3940_;
  assign new_n3956_ = new_n3955_ & new_n3926_;
  assign new_n3957_ = ~new_n3956_;
  assign new_n3958_ = new_n3957_ & new_n264_;
  assign new_n3959_ = ~new_n3958_;
  assign new_n3960_ = new_n1959_ & new_n267_;
  assign new_n3961_ = ~new_n3960_;
  assign new_n3962_ = new_n1974_ & new_n293_;
  assign new_n3963_ = ~new_n3962_;
  assign new_n3964_ = new_n3963_ & new_n3961_;
  assign new_n3965_ = new_n2021_ & new_n318_;
  assign new_n3966_ = ~new_n3965_;
  assign new_n3967_ = new_n1967_ & new_n342_;
  assign new_n3968_ = ~new_n3967_;
  assign new_n3969_ = new_n3968_ & new_n3966_;
  assign new_n3970_ = new_n3969_ & new_n3964_;
  assign new_n3971_ = ~new_n3970_;
  assign new_n3972_ = new_n3971_ & new_n669_;
  assign new_n3973_ = ~new_n3972_;
  assign new_n3974_ = new_n1817_ & new_n267_;
  assign new_n3975_ = ~new_n3974_;
  assign new_n3976_ = new_n1832_ & new_n293_;
  assign new_n3977_ = ~new_n3976_;
  assign new_n3978_ = new_n3977_ & new_n3975_;
  assign new_n3979_ = new_n1952_ & new_n318_;
  assign new_n3980_ = ~new_n3979_;
  assign new_n3981_ = new_n1825_ & new_n342_;
  assign new_n3982_ = ~new_n3981_;
  assign new_n3983_ = new_n3982_ & new_n3980_;
  assign new_n3984_ = new_n3983_ & new_n3978_;
  assign new_n3985_ = ~new_n3984_;
  assign new_n3986_ = new_n3985_ & new_n570_;
  assign new_n3987_ = ~new_n3986_;
  assign new_n3988_ = new_n3987_ & new_n3973_;
  assign new_n3989_ = new_n2028_ & new_n267_;
  assign new_n3990_ = ~new_n3989_;
  assign new_n3991_ = new_n2051_ & new_n293_;
  assign new_n3992_ = ~new_n3991_;
  assign new_n3993_ = new_n3992_ & new_n3990_;
  assign new_n3994_ = new_n2063_ & new_n318_;
  assign new_n3995_ = ~new_n3994_;
  assign new_n3996_ = new_n2040_ & new_n342_;
  assign new_n3997_ = ~new_n3996_;
  assign new_n3998_ = new_n3997_ & new_n3995_;
  assign new_n3999_ = new_n3998_ & new_n3993_;
  assign new_n4000_ = ~new_n3999_;
  assign new_n4001_ = new_n4000_ & new_n469_;
  assign new_n4002_ = ~new_n4001_;
  assign new_n4003_ = new_n2070_ & new_n267_;
  assign new_n4004_ = ~new_n4003_;
  assign new_n4005_ = new_n2085_ & new_n293_;
  assign new_n4006_ = ~new_n4005_;
  assign new_n4007_ = new_n4006_ & new_n4004_;
  assign new_n4008_ = new_n1986_ & new_n318_;
  assign new_n4009_ = ~new_n4008_;
  assign new_n4010_ = new_n2078_ & new_n342_;
  assign new_n4011_ = ~new_n4010_;
  assign new_n4012_ = new_n4011_ & new_n4009_;
  assign new_n4013_ = new_n4012_ & new_n4007_;
  assign new_n4014_ = ~new_n4013_;
  assign new_n4015_ = new_n4014_ & new_n369_;
  assign new_n4016_ = ~new_n4015_;
  assign new_n4017_ = new_n4016_ & new_n4002_;
  assign new_n4018_ = new_n4017_ & new_n3988_;
  assign new_n4019_ = ~new_n4018_;
  assign new_n4020_ = new_n4019_ & shift6;
  assign new_n4021_ = ~new_n4020_;
  assign new_n4022_ = new_n4021_ & new_n3959_;
  assign ores14 = ~new_n4022_;
  assign new_n4024_ = new_n2193_ & new_n267_;
  assign new_n4025_ = ~new_n4024_;
  assign new_n4026_ = new_n2224_ & new_n293_;
  assign new_n4027_ = ~new_n4026_;
  assign new_n4028_ = new_n4027_ & new_n4025_;
  assign new_n4029_ = new_n2311_ & new_n318_;
  assign new_n4030_ = ~new_n4029_;
  assign new_n4031_ = new_n2209_ & new_n342_;
  assign new_n4032_ = ~new_n4031_;
  assign new_n4033_ = new_n4032_ & new_n4030_;
  assign new_n4034_ = new_n4033_ & new_n4028_;
  assign new_n4035_ = ~new_n4034_;
  assign new_n4036_ = new_n4035_ & new_n369_;
  assign new_n4037_ = ~new_n4036_;
  assign new_n4038_ = new_n2127_ & new_n267_;
  assign new_n4039_ = ~new_n4038_;
  assign new_n4040_ = new_n2158_ & new_n293_;
  assign new_n4041_ = ~new_n4040_;
  assign new_n4042_ = new_n4041_ & new_n4039_;
  assign new_n4043_ = new_n2178_ & new_n318_;
  assign new_n4044_ = ~new_n4043_;
  assign new_n4045_ = new_n2143_ & new_n342_;
  assign new_n4046_ = ~new_n4045_;
  assign new_n4047_ = new_n4046_ & new_n4044_;
  assign new_n4048_ = new_n4047_ & new_n4042_;
  assign new_n4049_ = ~new_n4048_;
  assign new_n4050_ = new_n4049_ & new_n469_;
  assign new_n4051_ = ~new_n4050_;
  assign new_n4052_ = new_n4051_ & new_n4037_;
  assign new_n4053_ = new_n2526_ & new_n267_;
  assign new_n4054_ = ~new_n4053_;
  assign new_n4055_ = new_n2557_ & new_n293_;
  assign new_n4056_ = ~new_n4055_;
  assign new_n4057_ = new_n4056_ & new_n4054_;
  assign new_n4058_ = new_n2245_ & new_n318_;
  assign new_n4059_ = ~new_n4058_;
  assign new_n4060_ = new_n2542_ & new_n342_;
  assign new_n4061_ = ~new_n4060_;
  assign new_n4062_ = new_n4061_ & new_n4059_;
  assign new_n4063_ = new_n4062_ & new_n4057_;
  assign new_n4064_ = ~new_n4063_;
  assign new_n4065_ = new_n4064_ & new_n570_;
  assign new_n4066_ = ~new_n4065_;
  assign new_n4067_ = new_n2260_ & new_n267_;
  assign new_n4068_ = ~new_n4067_;
  assign new_n4069_ = new_n2291_ & new_n293_;
  assign new_n4070_ = ~new_n4069_;
  assign new_n4071_ = new_n4070_ & new_n4068_;
  assign new_n4072_ = new_n2112_ & new_n318_;
  assign new_n4073_ = ~new_n4072_;
  assign new_n4074_ = new_n2276_ & new_n342_;
  assign new_n4075_ = ~new_n4074_;
  assign new_n4076_ = new_n4075_ & new_n4073_;
  assign new_n4077_ = new_n4076_ & new_n4071_;
  assign new_n4078_ = ~new_n4077_;
  assign new_n4079_ = new_n4078_ & new_n669_;
  assign new_n4080_ = ~new_n4079_;
  assign new_n4081_ = new_n4080_ & new_n4066_;
  assign new_n4082_ = new_n4081_ & new_n4052_;
  assign new_n4083_ = ~new_n4082_;
  assign new_n4084_ = new_n4083_ & new_n264_;
  assign new_n4085_ = ~new_n4084_;
  assign new_n4086_ = new_n2397_ & new_n267_;
  assign new_n4087_ = ~new_n4086_;
  assign new_n4088_ = new_n2428_ & new_n293_;
  assign new_n4089_ = ~new_n4088_;
  assign new_n4090_ = new_n4089_ & new_n4087_;
  assign new_n4091_ = new_n2448_ & new_n318_;
  assign new_n4092_ = ~new_n4091_;
  assign new_n4093_ = new_n2413_ & new_n342_;
  assign new_n4094_ = ~new_n4093_;
  assign new_n4095_ = new_n4094_ & new_n4092_;
  assign new_n4096_ = new_n4095_ & new_n4090_;
  assign new_n4097_ = ~new_n4096_;
  assign new_n4098_ = new_n4097_ & new_n669_;
  assign new_n4099_ = ~new_n4098_;
  assign new_n4100_ = new_n2326_ & new_n267_;
  assign new_n4101_ = ~new_n4100_;
  assign new_n4102_ = new_n2357_ & new_n293_;
  assign new_n4103_ = ~new_n4102_;
  assign new_n4104_ = new_n4103_ & new_n4101_;
  assign new_n4105_ = new_n2382_ & new_n318_;
  assign new_n4106_ = ~new_n4105_;
  assign new_n4107_ = new_n2342_ & new_n342_;
  assign new_n4108_ = ~new_n4107_;
  assign new_n4109_ = new_n4108_ & new_n4106_;
  assign new_n4110_ = new_n4109_ & new_n4104_;
  assign new_n4111_ = ~new_n4110_;
  assign new_n4112_ = new_n4111_ & new_n570_;
  assign new_n4113_ = ~new_n4112_;
  assign new_n4114_ = new_n4113_ & new_n4099_;
  assign new_n4115_ = new_n2459_ & new_n267_;
  assign new_n4116_ = ~new_n4115_;
  assign new_n4117_ = new_n2490_ & new_n293_;
  assign new_n4118_ = ~new_n4117_;
  assign new_n4119_ = new_n4118_ & new_n4116_;
  assign new_n4120_ = new_n2577_ & new_n318_;
  assign new_n4121_ = ~new_n4120_;
  assign new_n4122_ = new_n2475_ & new_n342_;
  assign new_n4123_ = ~new_n4122_;
  assign new_n4124_ = new_n4123_ & new_n4121_;
  assign new_n4125_ = new_n4124_ & new_n4119_;
  assign new_n4126_ = ~new_n4125_;
  assign new_n4127_ = new_n4126_ & new_n469_;
  assign new_n4128_ = ~new_n4127_;
  assign new_n4129_ = new_n2592_ & new_n267_;
  assign new_n4130_ = ~new_n4129_;
  assign new_n4131_ = new_n2623_ & new_n293_;
  assign new_n4132_ = ~new_n4131_;
  assign new_n4133_ = new_n4132_ & new_n4130_;
  assign new_n4134_ = new_n2511_ & new_n318_;
  assign new_n4135_ = ~new_n4134_;
  assign new_n4136_ = new_n2608_ & new_n342_;
  assign new_n4137_ = ~new_n4136_;
  assign new_n4138_ = new_n4137_ & new_n4135_;
  assign new_n4139_ = new_n4138_ & new_n4133_;
  assign new_n4140_ = ~new_n4139_;
  assign new_n4141_ = new_n4140_ & new_n369_;
  assign new_n4142_ = ~new_n4141_;
  assign new_n4143_ = new_n4142_ & new_n4128_;
  assign new_n4144_ = new_n4143_ & new_n4114_;
  assign new_n4145_ = ~new_n4144_;
  assign new_n4146_ = new_n4145_ & shift6;
  assign new_n4147_ = ~new_n4146_;
  assign new_n4148_ = new_n4147_ & new_n4085_;
  assign ores15 = ~new_n4148_;
  assign new_n4150_ = new_n467_ & new_n369_;
  assign new_n4151_ = ~new_n4150_;
  assign new_n4152_ = new_n668_ & new_n469_;
  assign new_n4153_ = ~new_n4152_;
  assign new_n4154_ = new_n4153_ & new_n4151_;
  assign new_n4155_ = new_n772_ & new_n570_;
  assign new_n4156_ = ~new_n4155_;
  assign new_n4157_ = new_n669_ & new_n568_;
  assign new_n4158_ = ~new_n4157_;
  assign new_n4159_ = new_n4158_ & new_n4156_;
  assign new_n4160_ = new_n4159_ & new_n4154_;
  assign new_n4161_ = ~new_n4160_;
  assign new_n4162_ = new_n4161_ & new_n264_;
  assign new_n4163_ = ~new_n4162_;
  assign new_n4164_ = new_n570_ & new_n368_;
  assign new_n4165_ = ~new_n4164_;
  assign new_n4166_ = new_n870_ & new_n369_;
  assign new_n4167_ = ~new_n4166_;
  assign new_n4168_ = new_n4167_ & new_n4165_;
  assign new_n4169_ = new_n969_ & new_n669_;
  assign new_n4170_ = ~new_n4169_;
  assign new_n4171_ = new_n1065_ & new_n469_;
  assign new_n4172_ = ~new_n4171_;
  assign new_n4173_ = new_n4172_ & new_n4170_;
  assign new_n4174_ = new_n4173_ & new_n4168_;
  assign new_n4175_ = ~new_n4174_;
  assign new_n4176_ = new_n4175_ & shift6;
  assign new_n4177_ = ~new_n4176_;
  assign new_n4178_ = new_n4177_ & new_n4163_;
  assign ores16 = ~new_n4178_;
  assign new_n4180_ = new_n1252_ & new_n369_;
  assign new_n4181_ = ~new_n4180_;
  assign new_n4182_ = new_n1433_ & new_n469_;
  assign new_n4183_ = ~new_n4182_;
  assign new_n4184_ = new_n4183_ & new_n4181_;
  assign new_n4185_ = new_n1618_ & new_n570_;
  assign new_n4186_ = ~new_n4185_;
  assign new_n4187_ = new_n1343_ & new_n669_;
  assign new_n4188_ = ~new_n4187_;
  assign new_n4189_ = new_n4188_ & new_n4186_;
  assign new_n4190_ = new_n4189_ & new_n4184_;
  assign new_n4191_ = ~new_n4190_;
  assign new_n4192_ = new_n4191_ & new_n264_;
  assign new_n4193_ = ~new_n4192_;
  assign new_n4194_ = new_n1528_ & new_n669_;
  assign new_n4195_ = ~new_n4194_;
  assign new_n4196_ = new_n1162_ & new_n570_;
  assign new_n4197_ = ~new_n4196_;
  assign new_n4198_ = new_n4197_ & new_n4195_;
  assign new_n4199_ = new_n1706_ & new_n469_;
  assign new_n4200_ = ~new_n4199_;
  assign new_n4201_ = new_n1796_ & new_n369_;
  assign new_n4202_ = ~new_n4201_;
  assign new_n4203_ = new_n4202_ & new_n4200_;
  assign new_n4204_ = new_n4203_ & new_n4198_;
  assign new_n4205_ = ~new_n4204_;
  assign new_n4206_ = new_n4205_ & shift6;
  assign new_n4207_ = ~new_n4206_;
  assign new_n4208_ = new_n4207_ & new_n4193_;
  assign ores17 = ~new_n4208_;
  assign new_n4210_ = new_n1871_ & new_n369_;
  assign new_n4211_ = ~new_n4210_;
  assign new_n4212_ = new_n1940_ & new_n469_;
  assign new_n4213_ = ~new_n4212_;
  assign new_n4214_ = new_n4213_ & new_n4211_;
  assign new_n4215_ = new_n2013_ & new_n570_;
  assign new_n4216_ = ~new_n4215_;
  assign new_n4217_ = new_n1906_ & new_n669_;
  assign new_n4218_ = ~new_n4217_;
  assign new_n4219_ = new_n4218_ & new_n4216_;
  assign new_n4220_ = new_n4219_ & new_n4214_;
  assign new_n4221_ = ~new_n4220_;
  assign new_n4222_ = new_n4221_ & new_n264_;
  assign new_n4223_ = ~new_n4222_;
  assign new_n4224_ = new_n1979_ & new_n669_;
  assign new_n4225_ = ~new_n4224_;
  assign new_n4226_ = new_n1837_ & new_n570_;
  assign new_n4227_ = ~new_n4226_;
  assign new_n4228_ = new_n4227_ & new_n4225_;
  assign new_n4229_ = new_n2056_ & new_n469_;
  assign new_n4230_ = ~new_n4229_;
  assign new_n4231_ = new_n2090_ & new_n369_;
  assign new_n4232_ = ~new_n4231_;
  assign new_n4233_ = new_n4232_ & new_n4230_;
  assign new_n4234_ = new_n4233_ & new_n4228_;
  assign new_n4235_ = ~new_n4234_;
  assign new_n4236_ = new_n4235_ & shift6;
  assign new_n4237_ = ~new_n4236_;
  assign new_n4238_ = new_n4237_ & new_n4223_;
  assign ores18 = ~new_n4238_;
  assign new_n4240_ = new_n2163_ & new_n469_;
  assign new_n4241_ = ~new_n4240_;
  assign new_n4242_ = new_n2229_ & new_n369_;
  assign new_n4243_ = ~new_n4242_;
  assign new_n4244_ = new_n4243_ & new_n4241_;
  assign new_n4245_ = new_n2296_ & new_n669_;
  assign new_n4246_ = ~new_n4245_;
  assign new_n4247_ = new_n2562_ & new_n570_;
  assign new_n4248_ = ~new_n4247_;
  assign new_n4249_ = new_n4248_ & new_n4246_;
  assign new_n4250_ = new_n4249_ & new_n4244_;
  assign new_n4251_ = ~new_n4250_;
  assign new_n4252_ = new_n4251_ & new_n264_;
  assign new_n4253_ = ~new_n4252_;
  assign new_n4254_ = new_n2433_ & new_n669_;
  assign new_n4255_ = ~new_n4254_;
  assign new_n4256_ = new_n2362_ & new_n570_;
  assign new_n4257_ = ~new_n4256_;
  assign new_n4258_ = new_n4257_ & new_n4255_;
  assign new_n4259_ = new_n2628_ & new_n369_;
  assign new_n4260_ = ~new_n4259_;
  assign new_n4261_ = new_n2495_ & new_n469_;
  assign new_n4262_ = ~new_n4261_;
  assign new_n4263_ = new_n4262_ & new_n4260_;
  assign new_n4264_ = new_n4263_ & new_n4258_;
  assign new_n4265_ = ~new_n4264_;
  assign new_n4266_ = new_n4265_ & shift6;
  assign new_n4267_ = ~new_n4266_;
  assign new_n4268_ = new_n4267_ & new_n4253_;
  assign ores19 = ~new_n4268_;
  assign new_n4270_ = new_n2663_ & new_n369_;
  assign new_n4271_ = ~new_n4270_;
  assign new_n4272_ = new_n2692_ & new_n469_;
  assign new_n4273_ = ~new_n4272_;
  assign new_n4274_ = new_n4273_ & new_n4271_;
  assign new_n4275_ = new_n2754_ & new_n570_;
  assign new_n4276_ = ~new_n4275_;
  assign new_n4277_ = new_n2678_ & new_n669_;
  assign new_n4278_ = ~new_n4277_;
  assign new_n4279_ = new_n4278_ & new_n4276_;
  assign new_n4280_ = new_n4279_ & new_n4274_;
  assign new_n4281_ = ~new_n4280_;
  assign new_n4282_ = new_n4281_ & new_n264_;
  assign new_n4283_ = ~new_n4282_;
  assign new_n4284_ = new_n2649_ & new_n570_;
  assign new_n4285_ = ~new_n4284_;
  assign new_n4286_ = new_n2711_ & new_n469_;
  assign new_n4287_ = ~new_n4286_;
  assign new_n4288_ = new_n4287_ & new_n4285_;
  assign new_n4289_ = new_n2740_ & new_n369_;
  assign new_n4290_ = ~new_n4289_;
  assign new_n4291_ = new_n2725_ & new_n669_;
  assign new_n4292_ = ~new_n4291_;
  assign new_n4293_ = new_n4292_ & new_n4290_;
  assign new_n4294_ = new_n4293_ & new_n4288_;
  assign new_n4295_ = ~new_n4294_;
  assign new_n4296_ = new_n4295_ & shift6;
  assign new_n4297_ = ~new_n4296_;
  assign new_n4298_ = new_n4297_ & new_n4283_;
  assign ores20 = ~new_n4298_;
  assign new_n4300_ = new_n2789_ & new_n369_;
  assign new_n4301_ = ~new_n4300_;
  assign new_n4302_ = new_n2818_ & new_n469_;
  assign new_n4303_ = ~new_n4302_;
  assign new_n4304_ = new_n4303_ & new_n4301_;
  assign new_n4305_ = new_n2880_ & new_n570_;
  assign new_n4306_ = ~new_n4305_;
  assign new_n4307_ = new_n2804_ & new_n669_;
  assign new_n4308_ = ~new_n4307_;
  assign new_n4309_ = new_n4308_ & new_n4306_;
  assign new_n4310_ = new_n4309_ & new_n4304_;
  assign new_n4311_ = ~new_n4310_;
  assign new_n4312_ = new_n4311_ & new_n264_;
  assign new_n4313_ = ~new_n4312_;
  assign new_n4314_ = new_n2775_ & new_n570_;
  assign new_n4315_ = ~new_n4314_;
  assign new_n4316_ = new_n2837_ & new_n469_;
  assign new_n4317_ = ~new_n4316_;
  assign new_n4318_ = new_n4317_ & new_n4315_;
  assign new_n4319_ = new_n2866_ & new_n369_;
  assign new_n4320_ = ~new_n4319_;
  assign new_n4321_ = new_n2851_ & new_n669_;
  assign new_n4322_ = ~new_n4321_;
  assign new_n4323_ = new_n4322_ & new_n4320_;
  assign new_n4324_ = new_n4323_ & new_n4318_;
  assign new_n4325_ = ~new_n4324_;
  assign new_n4326_ = new_n4325_ & shift6;
  assign new_n4327_ = ~new_n4326_;
  assign new_n4328_ = new_n4327_ & new_n4313_;
  assign ores21 = ~new_n4328_;
  assign new_n4330_ = new_n2915_ & new_n369_;
  assign new_n4331_ = ~new_n4330_;
  assign new_n4332_ = new_n2944_ & new_n469_;
  assign new_n4333_ = ~new_n4332_;
  assign new_n4334_ = new_n4333_ & new_n4331_;
  assign new_n4335_ = new_n3006_ & new_n570_;
  assign new_n4336_ = ~new_n4335_;
  assign new_n4337_ = new_n2930_ & new_n669_;
  assign new_n4338_ = ~new_n4337_;
  assign new_n4339_ = new_n4338_ & new_n4336_;
  assign new_n4340_ = new_n4339_ & new_n4334_;
  assign new_n4341_ = ~new_n4340_;
  assign new_n4342_ = new_n4341_ & new_n264_;
  assign new_n4343_ = ~new_n4342_;
  assign new_n4344_ = new_n2901_ & new_n570_;
  assign new_n4345_ = ~new_n4344_;
  assign new_n4346_ = new_n2963_ & new_n469_;
  assign new_n4347_ = ~new_n4346_;
  assign new_n4348_ = new_n4347_ & new_n4345_;
  assign new_n4349_ = new_n2992_ & new_n369_;
  assign new_n4350_ = ~new_n4349_;
  assign new_n4351_ = new_n2977_ & new_n669_;
  assign new_n4352_ = ~new_n4351_;
  assign new_n4353_ = new_n4352_ & new_n4350_;
  assign new_n4354_ = new_n4353_ & new_n4348_;
  assign new_n4355_ = ~new_n4354_;
  assign new_n4356_ = new_n4355_ & shift6;
  assign new_n4357_ = ~new_n4356_;
  assign new_n4358_ = new_n4357_ & new_n4343_;
  assign ores22 = ~new_n4358_;
  assign new_n4360_ = new_n3041_ & new_n369_;
  assign new_n4361_ = ~new_n4360_;
  assign new_n4362_ = new_n3132_ & new_n570_;
  assign new_n4363_ = ~new_n4362_;
  assign new_n4364_ = new_n4363_ & new_n4361_;
  assign new_n4365_ = new_n3056_ & new_n669_;
  assign new_n4366_ = ~new_n4365_;
  assign new_n4367_ = new_n3070_ & new_n469_;
  assign new_n4368_ = ~new_n4367_;
  assign new_n4369_ = new_n4368_ & new_n4366_;
  assign new_n4370_ = new_n4369_ & new_n4364_;
  assign new_n4371_ = ~new_n4370_;
  assign new_n4372_ = new_n4371_ & new_n264_;
  assign new_n4373_ = ~new_n4372_;
  assign new_n4374_ = new_n3089_ & new_n469_;
  assign new_n4375_ = ~new_n4374_;
  assign new_n4376_ = new_n3103_ & new_n669_;
  assign new_n4377_ = ~new_n4376_;
  assign new_n4378_ = new_n4377_ & new_n4375_;
  assign new_n4379_ = new_n3118_ & new_n369_;
  assign new_n4380_ = ~new_n4379_;
  assign new_n4381_ = new_n3027_ & new_n570_;
  assign new_n4382_ = ~new_n4381_;
  assign new_n4383_ = new_n4382_ & new_n4380_;
  assign new_n4384_ = new_n4383_ & new_n4378_;
  assign new_n4385_ = ~new_n4384_;
  assign new_n4386_ = new_n4385_ & shift6;
  assign new_n4387_ = ~new_n4386_;
  assign new_n4388_ = new_n4387_ & new_n4373_;
  assign ores23 = ~new_n4388_;
  assign new_n4390_ = new_n3167_ & new_n369_;
  assign new_n4391_ = ~new_n4390_;
  assign new_n4392_ = new_n3258_ & new_n570_;
  assign new_n4393_ = ~new_n4392_;
  assign new_n4394_ = new_n4393_ & new_n4391_;
  assign new_n4395_ = new_n3182_ & new_n669_;
  assign new_n4396_ = ~new_n4395_;
  assign new_n4397_ = new_n3196_ & new_n469_;
  assign new_n4398_ = ~new_n4397_;
  assign new_n4399_ = new_n4398_ & new_n4396_;
  assign new_n4400_ = new_n4399_ & new_n4394_;
  assign new_n4401_ = ~new_n4400_;
  assign new_n4402_ = new_n4401_ & new_n264_;
  assign new_n4403_ = ~new_n4402_;
  assign new_n4404_ = new_n3215_ & new_n469_;
  assign new_n4405_ = ~new_n4404_;
  assign new_n4406_ = new_n3229_ & new_n669_;
  assign new_n4407_ = ~new_n4406_;
  assign new_n4408_ = new_n4407_ & new_n4405_;
  assign new_n4409_ = new_n3244_ & new_n369_;
  assign new_n4410_ = ~new_n4409_;
  assign new_n4411_ = new_n3153_ & new_n570_;
  assign new_n4412_ = ~new_n4411_;
  assign new_n4413_ = new_n4412_ & new_n4410_;
  assign new_n4414_ = new_n4413_ & new_n4408_;
  assign new_n4415_ = ~new_n4414_;
  assign new_n4416_ = new_n4415_ & shift6;
  assign new_n4417_ = ~new_n4416_;
  assign new_n4418_ = new_n4417_ & new_n4403_;
  assign ores24 = ~new_n4418_;
  assign new_n4420_ = new_n3293_ & new_n369_;
  assign new_n4421_ = ~new_n4420_;
  assign new_n4422_ = new_n3384_ & new_n570_;
  assign new_n4423_ = ~new_n4422_;
  assign new_n4424_ = new_n4423_ & new_n4421_;
  assign new_n4425_ = new_n3308_ & new_n669_;
  assign new_n4426_ = ~new_n4425_;
  assign new_n4427_ = new_n3322_ & new_n469_;
  assign new_n4428_ = ~new_n4427_;
  assign new_n4429_ = new_n4428_ & new_n4426_;
  assign new_n4430_ = new_n4429_ & new_n4424_;
  assign new_n4431_ = ~new_n4430_;
  assign new_n4432_ = new_n4431_ & new_n264_;
  assign new_n4433_ = ~new_n4432_;
  assign new_n4434_ = new_n3341_ & new_n469_;
  assign new_n4435_ = ~new_n4434_;
  assign new_n4436_ = new_n3355_ & new_n669_;
  assign new_n4437_ = ~new_n4436_;
  assign new_n4438_ = new_n4437_ & new_n4435_;
  assign new_n4439_ = new_n3370_ & new_n369_;
  assign new_n4440_ = ~new_n4439_;
  assign new_n4441_ = new_n3279_ & new_n570_;
  assign new_n4442_ = ~new_n4441_;
  assign new_n4443_ = new_n4442_ & new_n4440_;
  assign new_n4444_ = new_n4443_ & new_n4438_;
  assign new_n4445_ = ~new_n4444_;
  assign new_n4446_ = new_n4445_ & shift6;
  assign new_n4447_ = ~new_n4446_;
  assign new_n4448_ = new_n4447_ & new_n4433_;
  assign ores25 = ~new_n4448_;
  assign new_n4450_ = new_n3419_ & new_n369_;
  assign new_n4451_ = ~new_n4450_;
  assign new_n4452_ = new_n3448_ & new_n469_;
  assign new_n4453_ = ~new_n4452_;
  assign new_n4454_ = new_n4453_ & new_n4451_;
  assign new_n4455_ = new_n3510_ & new_n570_;
  assign new_n4456_ = ~new_n4455_;
  assign new_n4457_ = new_n3434_ & new_n669_;
  assign new_n4458_ = ~new_n4457_;
  assign new_n4459_ = new_n4458_ & new_n4456_;
  assign new_n4460_ = new_n4459_ & new_n4454_;
  assign new_n4461_ = ~new_n4460_;
  assign new_n4462_ = new_n4461_ & new_n264_;
  assign new_n4463_ = ~new_n4462_;
  assign new_n4464_ = new_n3467_ & new_n469_;
  assign new_n4465_ = ~new_n4464_;
  assign new_n4466_ = new_n3481_ & new_n669_;
  assign new_n4467_ = ~new_n4466_;
  assign new_n4468_ = new_n4467_ & new_n4465_;
  assign new_n4469_ = new_n3496_ & new_n369_;
  assign new_n4470_ = ~new_n4469_;
  assign new_n4471_ = new_n3405_ & new_n570_;
  assign new_n4472_ = ~new_n4471_;
  assign new_n4473_ = new_n4472_ & new_n4470_;
  assign new_n4474_ = new_n4473_ & new_n4468_;
  assign new_n4475_ = ~new_n4474_;
  assign new_n4476_ = new_n4475_ & shift6;
  assign new_n4477_ = ~new_n4476_;
  assign new_n4478_ = new_n4477_ & new_n4463_;
  assign ores26 = ~new_n4478_;
  assign new_n4480_ = new_n3545_ & new_n369_;
  assign new_n4481_ = ~new_n4480_;
  assign new_n4482_ = new_n3574_ & new_n469_;
  assign new_n4483_ = ~new_n4482_;
  assign new_n4484_ = new_n4483_ & new_n4481_;
  assign new_n4485_ = new_n3636_ & new_n570_;
  assign new_n4486_ = ~new_n4485_;
  assign new_n4487_ = new_n3560_ & new_n669_;
  assign new_n4488_ = ~new_n4487_;
  assign new_n4489_ = new_n4488_ & new_n4486_;
  assign new_n4490_ = new_n4489_ & new_n4484_;
  assign new_n4491_ = ~new_n4490_;
  assign new_n4492_ = new_n4491_ & new_n264_;
  assign new_n4493_ = ~new_n4492_;
  assign new_n4494_ = new_n3593_ & new_n469_;
  assign new_n4495_ = ~new_n4494_;
  assign new_n4496_ = new_n3607_ & new_n669_;
  assign new_n4497_ = ~new_n4496_;
  assign new_n4498_ = new_n4497_ & new_n4495_;
  assign new_n4499_ = new_n3622_ & new_n369_;
  assign new_n4500_ = ~new_n4499_;
  assign new_n4501_ = new_n3531_ & new_n570_;
  assign new_n4502_ = ~new_n4501_;
  assign new_n4503_ = new_n4502_ & new_n4500_;
  assign new_n4504_ = new_n4503_ & new_n4498_;
  assign new_n4505_ = ~new_n4504_;
  assign new_n4506_ = new_n4505_ & shift6;
  assign new_n4507_ = ~new_n4506_;
  assign new_n4508_ = new_n4507_ & new_n4493_;
  assign ores27 = ~new_n4508_;
  assign new_n4510_ = new_n3671_ & new_n369_;
  assign new_n4511_ = ~new_n4510_;
  assign new_n4512_ = new_n3700_ & new_n469_;
  assign new_n4513_ = ~new_n4512_;
  assign new_n4514_ = new_n4513_ & new_n4511_;
  assign new_n4515_ = new_n3762_ & new_n570_;
  assign new_n4516_ = ~new_n4515_;
  assign new_n4517_ = new_n3686_ & new_n669_;
  assign new_n4518_ = ~new_n4517_;
  assign new_n4519_ = new_n4518_ & new_n4516_;
  assign new_n4520_ = new_n4519_ & new_n4514_;
  assign new_n4521_ = ~new_n4520_;
  assign new_n4522_ = new_n4521_ & new_n264_;
  assign new_n4523_ = ~new_n4522_;
  assign new_n4524_ = new_n3719_ & new_n469_;
  assign new_n4525_ = ~new_n4524_;
  assign new_n4526_ = new_n3733_ & new_n669_;
  assign new_n4527_ = ~new_n4526_;
  assign new_n4528_ = new_n4527_ & new_n4525_;
  assign new_n4529_ = new_n3748_ & new_n369_;
  assign new_n4530_ = ~new_n4529_;
  assign new_n4531_ = new_n3657_ & new_n570_;
  assign new_n4532_ = ~new_n4531_;
  assign new_n4533_ = new_n4532_ & new_n4530_;
  assign new_n4534_ = new_n4533_ & new_n4528_;
  assign new_n4535_ = ~new_n4534_;
  assign new_n4536_ = new_n4535_ & shift6;
  assign new_n4537_ = ~new_n4536_;
  assign new_n4538_ = new_n4537_ & new_n4523_;
  assign ores28 = ~new_n4538_;
  assign new_n4540_ = new_n3797_ & new_n369_;
  assign new_n4541_ = ~new_n4540_;
  assign new_n4542_ = new_n3826_ & new_n469_;
  assign new_n4543_ = ~new_n4542_;
  assign new_n4544_ = new_n4543_ & new_n4541_;
  assign new_n4545_ = new_n3888_ & new_n570_;
  assign new_n4546_ = ~new_n4545_;
  assign new_n4547_ = new_n3812_ & new_n669_;
  assign new_n4548_ = ~new_n4547_;
  assign new_n4549_ = new_n4548_ & new_n4546_;
  assign new_n4550_ = new_n4549_ & new_n4544_;
  assign new_n4551_ = ~new_n4550_;
  assign new_n4552_ = new_n4551_ & new_n264_;
  assign new_n4553_ = ~new_n4552_;
  assign new_n4554_ = new_n3845_ & new_n469_;
  assign new_n4555_ = ~new_n4554_;
  assign new_n4556_ = new_n3859_ & new_n669_;
  assign new_n4557_ = ~new_n4556_;
  assign new_n4558_ = new_n4557_ & new_n4555_;
  assign new_n4559_ = new_n3874_ & new_n369_;
  assign new_n4560_ = ~new_n4559_;
  assign new_n4561_ = new_n3783_ & new_n570_;
  assign new_n4562_ = ~new_n4561_;
  assign new_n4563_ = new_n4562_ & new_n4560_;
  assign new_n4564_ = new_n4563_ & new_n4558_;
  assign new_n4565_ = ~new_n4564_;
  assign new_n4566_ = new_n4565_ & shift6;
  assign new_n4567_ = ~new_n4566_;
  assign new_n4568_ = new_n4567_ & new_n4553_;
  assign ores29 = ~new_n4568_;
  assign new_n4570_ = new_n3923_ & new_n369_;
  assign new_n4571_ = ~new_n4570_;
  assign new_n4572_ = new_n3952_ & new_n469_;
  assign new_n4573_ = ~new_n4572_;
  assign new_n4574_ = new_n4573_ & new_n4571_;
  assign new_n4575_ = new_n4014_ & new_n570_;
  assign new_n4576_ = ~new_n4575_;
  assign new_n4577_ = new_n3938_ & new_n669_;
  assign new_n4578_ = ~new_n4577_;
  assign new_n4579_ = new_n4578_ & new_n4576_;
  assign new_n4580_ = new_n4579_ & new_n4574_;
  assign new_n4581_ = ~new_n4580_;
  assign new_n4582_ = new_n4581_ & new_n264_;
  assign new_n4583_ = ~new_n4582_;
  assign new_n4584_ = new_n3971_ & new_n469_;
  assign new_n4585_ = ~new_n4584_;
  assign new_n4586_ = new_n3985_ & new_n669_;
  assign new_n4587_ = ~new_n4586_;
  assign new_n4588_ = new_n4587_ & new_n4585_;
  assign new_n4589_ = new_n4000_ & new_n369_;
  assign new_n4590_ = ~new_n4589_;
  assign new_n4591_ = new_n3909_ & new_n570_;
  assign new_n4592_ = ~new_n4591_;
  assign new_n4593_ = new_n4592_ & new_n4590_;
  assign new_n4594_ = new_n4593_ & new_n4588_;
  assign new_n4595_ = ~new_n4594_;
  assign new_n4596_ = new_n4595_ & shift6;
  assign new_n4597_ = ~new_n4596_;
  assign new_n4598_ = new_n4597_ & new_n4583_;
  assign ores30 = ~new_n4598_;
  assign new_n4600_ = new_n4049_ & new_n369_;
  assign new_n4601_ = ~new_n4600_;
  assign new_n4602_ = new_n4078_ & new_n469_;
  assign new_n4603_ = ~new_n4602_;
  assign new_n4604_ = new_n4603_ & new_n4601_;
  assign new_n4605_ = new_n4140_ & new_n570_;
  assign new_n4606_ = ~new_n4605_;
  assign new_n4607_ = new_n4064_ & new_n669_;
  assign new_n4608_ = ~new_n4607_;
  assign new_n4609_ = new_n4608_ & new_n4606_;
  assign new_n4610_ = new_n4609_ & new_n4604_;
  assign new_n4611_ = ~new_n4610_;
  assign new_n4612_ = new_n4611_ & new_n264_;
  assign new_n4613_ = ~new_n4612_;
  assign new_n4614_ = new_n4097_ & new_n469_;
  assign new_n4615_ = ~new_n4614_;
  assign new_n4616_ = new_n4111_ & new_n669_;
  assign new_n4617_ = ~new_n4616_;
  assign new_n4618_ = new_n4617_ & new_n4615_;
  assign new_n4619_ = new_n4126_ & new_n369_;
  assign new_n4620_ = ~new_n4619_;
  assign new_n4621_ = new_n4035_ & new_n570_;
  assign new_n4622_ = ~new_n4621_;
  assign new_n4623_ = new_n4622_ & new_n4620_;
  assign new_n4624_ = new_n4623_ & new_n4618_;
  assign new_n4625_ = ~new_n4624_;
  assign new_n4626_ = new_n4625_ & shift6;
  assign new_n4627_ = ~new_n4626_;
  assign new_n4628_ = new_n4627_ & new_n4613_;
  assign ores31 = ~new_n4628_;
  assign new_n4630_ = new_n668_ & new_n369_;
  assign new_n4631_ = ~new_n4630_;
  assign new_n4632_ = new_n568_ & new_n469_;
  assign new_n4633_ = ~new_n4632_;
  assign new_n4634_ = new_n4633_ & new_n4631_;
  assign new_n4635_ = new_n870_ & new_n570_;
  assign new_n4636_ = ~new_n4635_;
  assign new_n4637_ = new_n772_ & new_n669_;
  assign new_n4638_ = ~new_n4637_;
  assign new_n4639_ = new_n4638_ & new_n4636_;
  assign new_n4640_ = new_n4639_ & new_n4634_;
  assign new_n4641_ = ~new_n4640_;
  assign new_n4642_ = new_n4641_ & new_n264_;
  assign new_n4643_ = ~new_n4642_;
  assign new_n4644_ = new_n669_ & new_n368_;
  assign new_n4645_ = ~new_n4644_;
  assign new_n4646_ = new_n570_ & new_n467_;
  assign new_n4647_ = ~new_n4646_;
  assign new_n4648_ = new_n4647_ & new_n4645_;
  assign new_n4649_ = new_n969_ & new_n469_;
  assign new_n4650_ = ~new_n4649_;
  assign new_n4651_ = new_n1065_ & new_n369_;
  assign new_n4652_ = ~new_n4651_;
  assign new_n4653_ = new_n4652_ & new_n4650_;
  assign new_n4654_ = new_n4653_ & new_n4648_;
  assign new_n4655_ = ~new_n4654_;
  assign new_n4656_ = new_n4655_ & shift6;
  assign new_n4657_ = ~new_n4656_;
  assign new_n4658_ = new_n4657_ & new_n4643_;
  assign ores32 = ~new_n4658_;
  assign new_n4660_ = new_n1433_ & new_n369_;
  assign new_n4661_ = ~new_n4660_;
  assign new_n4662_ = new_n1343_ & new_n469_;
  assign new_n4663_ = ~new_n4662_;
  assign new_n4664_ = new_n4663_ & new_n4661_;
  assign new_n4665_ = new_n1796_ & new_n570_;
  assign new_n4666_ = ~new_n4665_;
  assign new_n4667_ = new_n1618_ & new_n669_;
  assign new_n4668_ = ~new_n4667_;
  assign new_n4669_ = new_n4668_ & new_n4666_;
  assign new_n4670_ = new_n4669_ & new_n4664_;
  assign new_n4671_ = ~new_n4670_;
  assign new_n4672_ = new_n4671_ & new_n264_;
  assign new_n4673_ = ~new_n4672_;
  assign new_n4674_ = new_n1528_ & new_n469_;
  assign new_n4675_ = ~new_n4674_;
  assign new_n4676_ = new_n1162_ & new_n669_;
  assign new_n4677_ = ~new_n4676_;
  assign new_n4678_ = new_n4677_ & new_n4675_;
  assign new_n4679_ = new_n1706_ & new_n369_;
  assign new_n4680_ = ~new_n4679_;
  assign new_n4681_ = new_n1252_ & new_n570_;
  assign new_n4682_ = ~new_n4681_;
  assign new_n4683_ = new_n4682_ & new_n4680_;
  assign new_n4684_ = new_n4683_ & new_n4678_;
  assign new_n4685_ = ~new_n4684_;
  assign new_n4686_ = new_n4685_ & shift6;
  assign new_n4687_ = ~new_n4686_;
  assign new_n4688_ = new_n4687_ & new_n4673_;
  assign ores33 = ~new_n4688_;
  assign new_n4690_ = new_n1940_ & new_n369_;
  assign new_n4691_ = ~new_n4690_;
  assign new_n4692_ = new_n1906_ & new_n469_;
  assign new_n4693_ = ~new_n4692_;
  assign new_n4694_ = new_n4693_ & new_n4691_;
  assign new_n4695_ = new_n2090_ & new_n570_;
  assign new_n4696_ = ~new_n4695_;
  assign new_n4697_ = new_n2013_ & new_n669_;
  assign new_n4698_ = ~new_n4697_;
  assign new_n4699_ = new_n4698_ & new_n4696_;
  assign new_n4700_ = new_n4699_ & new_n4694_;
  assign new_n4701_ = ~new_n4700_;
  assign new_n4702_ = new_n4701_ & new_n264_;
  assign new_n4703_ = ~new_n4702_;
  assign new_n4704_ = new_n1979_ & new_n469_;
  assign new_n4705_ = ~new_n4704_;
  assign new_n4706_ = new_n1837_ & new_n669_;
  assign new_n4707_ = ~new_n4706_;
  assign new_n4708_ = new_n4707_ & new_n4705_;
  assign new_n4709_ = new_n2056_ & new_n369_;
  assign new_n4710_ = ~new_n4709_;
  assign new_n4711_ = new_n1871_ & new_n570_;
  assign new_n4712_ = ~new_n4711_;
  assign new_n4713_ = new_n4712_ & new_n4710_;
  assign new_n4714_ = new_n4713_ & new_n4708_;
  assign new_n4715_ = ~new_n4714_;
  assign new_n4716_ = new_n4715_ & shift6;
  assign new_n4717_ = ~new_n4716_;
  assign new_n4718_ = new_n4717_ & new_n4703_;
  assign ores34 = ~new_n4718_;
  assign new_n4720_ = new_n2163_ & new_n369_;
  assign new_n4721_ = ~new_n4720_;
  assign new_n4722_ = new_n2628_ & new_n570_;
  assign new_n4723_ = ~new_n4722_;
  assign new_n4724_ = new_n4723_ & new_n4721_;
  assign new_n4725_ = new_n2296_ & new_n469_;
  assign new_n4726_ = ~new_n4725_;
  assign new_n4727_ = new_n2562_ & new_n669_;
  assign new_n4728_ = ~new_n4727_;
  assign new_n4729_ = new_n4728_ & new_n4726_;
  assign new_n4730_ = new_n4729_ & new_n4724_;
  assign new_n4731_ = ~new_n4730_;
  assign new_n4732_ = new_n4731_ & new_n264_;
  assign new_n4733_ = ~new_n4732_;
  assign new_n4734_ = new_n2433_ & new_n469_;
  assign new_n4735_ = ~new_n4734_;
  assign new_n4736_ = new_n2229_ & new_n570_;
  assign new_n4737_ = ~new_n4736_;
  assign new_n4738_ = new_n4737_ & new_n4735_;
  assign new_n4739_ = new_n2495_ & new_n369_;
  assign new_n4740_ = ~new_n4739_;
  assign new_n4741_ = new_n2362_ & new_n669_;
  assign new_n4742_ = ~new_n4741_;
  assign new_n4743_ = new_n4742_ & new_n4740_;
  assign new_n4744_ = new_n4743_ & new_n4738_;
  assign new_n4745_ = ~new_n4744_;
  assign new_n4746_ = new_n4745_ & shift6;
  assign new_n4747_ = ~new_n4746_;
  assign new_n4748_ = new_n4747_ & new_n4733_;
  assign ores35 = ~new_n4748_;
  assign new_n4750_ = new_n2692_ & new_n369_;
  assign new_n4751_ = ~new_n4750_;
  assign new_n4752_ = new_n2678_ & new_n469_;
  assign new_n4753_ = ~new_n4752_;
  assign new_n4754_ = new_n4753_ & new_n4751_;
  assign new_n4755_ = new_n2740_ & new_n570_;
  assign new_n4756_ = ~new_n4755_;
  assign new_n4757_ = new_n2754_ & new_n669_;
  assign new_n4758_ = ~new_n4757_;
  assign new_n4759_ = new_n4758_ & new_n4756_;
  assign new_n4760_ = new_n4759_ & new_n4754_;
  assign new_n4761_ = ~new_n4760_;
  assign new_n4762_ = new_n4761_ & new_n264_;
  assign new_n4763_ = ~new_n4762_;
  assign new_n4764_ = new_n2649_ & new_n669_;
  assign new_n4765_ = ~new_n4764_;
  assign new_n4766_ = new_n2663_ & new_n570_;
  assign new_n4767_ = ~new_n4766_;
  assign new_n4768_ = new_n4767_ & new_n4765_;
  assign new_n4769_ = new_n2725_ & new_n469_;
  assign new_n4770_ = ~new_n4769_;
  assign new_n4771_ = new_n2711_ & new_n369_;
  assign new_n4772_ = ~new_n4771_;
  assign new_n4773_ = new_n4772_ & new_n4770_;
  assign new_n4774_ = new_n4773_ & new_n4768_;
  assign new_n4775_ = ~new_n4774_;
  assign new_n4776_ = new_n4775_ & shift6;
  assign new_n4777_ = ~new_n4776_;
  assign new_n4778_ = new_n4777_ & new_n4763_;
  assign ores36 = ~new_n4778_;
  assign new_n4780_ = new_n2818_ & new_n369_;
  assign new_n4781_ = ~new_n4780_;
  assign new_n4782_ = new_n2804_ & new_n469_;
  assign new_n4783_ = ~new_n4782_;
  assign new_n4784_ = new_n4783_ & new_n4781_;
  assign new_n4785_ = new_n2866_ & new_n570_;
  assign new_n4786_ = ~new_n4785_;
  assign new_n4787_ = new_n2880_ & new_n669_;
  assign new_n4788_ = ~new_n4787_;
  assign new_n4789_ = new_n4788_ & new_n4786_;
  assign new_n4790_ = new_n4789_ & new_n4784_;
  assign new_n4791_ = ~new_n4790_;
  assign new_n4792_ = new_n4791_ & new_n264_;
  assign new_n4793_ = ~new_n4792_;
  assign new_n4794_ = new_n2775_ & new_n669_;
  assign new_n4795_ = ~new_n4794_;
  assign new_n4796_ = new_n2789_ & new_n570_;
  assign new_n4797_ = ~new_n4796_;
  assign new_n4798_ = new_n4797_ & new_n4795_;
  assign new_n4799_ = new_n2851_ & new_n469_;
  assign new_n4800_ = ~new_n4799_;
  assign new_n4801_ = new_n2837_ & new_n369_;
  assign new_n4802_ = ~new_n4801_;
  assign new_n4803_ = new_n4802_ & new_n4800_;
  assign new_n4804_ = new_n4803_ & new_n4798_;
  assign new_n4805_ = ~new_n4804_;
  assign new_n4806_ = new_n4805_ & shift6;
  assign new_n4807_ = ~new_n4806_;
  assign new_n4808_ = new_n4807_ & new_n4793_;
  assign ores37 = ~new_n4808_;
  assign new_n4810_ = new_n2944_ & new_n369_;
  assign new_n4811_ = ~new_n4810_;
  assign new_n4812_ = new_n2930_ & new_n469_;
  assign new_n4813_ = ~new_n4812_;
  assign new_n4814_ = new_n4813_ & new_n4811_;
  assign new_n4815_ = new_n2992_ & new_n570_;
  assign new_n4816_ = ~new_n4815_;
  assign new_n4817_ = new_n3006_ & new_n669_;
  assign new_n4818_ = ~new_n4817_;
  assign new_n4819_ = new_n4818_ & new_n4816_;
  assign new_n4820_ = new_n4819_ & new_n4814_;
  assign new_n4821_ = ~new_n4820_;
  assign new_n4822_ = new_n4821_ & new_n264_;
  assign new_n4823_ = ~new_n4822_;
  assign new_n4824_ = new_n2901_ & new_n669_;
  assign new_n4825_ = ~new_n4824_;
  assign new_n4826_ = new_n2915_ & new_n570_;
  assign new_n4827_ = ~new_n4826_;
  assign new_n4828_ = new_n4827_ & new_n4825_;
  assign new_n4829_ = new_n2977_ & new_n469_;
  assign new_n4830_ = ~new_n4829_;
  assign new_n4831_ = new_n2963_ & new_n369_;
  assign new_n4832_ = ~new_n4831_;
  assign new_n4833_ = new_n4832_ & new_n4830_;
  assign new_n4834_ = new_n4833_ & new_n4828_;
  assign new_n4835_ = ~new_n4834_;
  assign new_n4836_ = new_n4835_ & shift6;
  assign new_n4837_ = ~new_n4836_;
  assign new_n4838_ = new_n4837_ & new_n4823_;
  assign ores38 = ~new_n4838_;
  assign new_n4840_ = new_n3132_ & new_n669_;
  assign new_n4841_ = ~new_n4840_;
  assign new_n4842_ = new_n3118_ & new_n570_;
  assign new_n4843_ = ~new_n4842_;
  assign new_n4844_ = new_n4843_ & new_n4841_;
  assign new_n4845_ = new_n3056_ & new_n469_;
  assign new_n4846_ = ~new_n4845_;
  assign new_n4847_ = new_n3070_ & new_n369_;
  assign new_n4848_ = ~new_n4847_;
  assign new_n4849_ = new_n4848_ & new_n4846_;
  assign new_n4850_ = new_n4849_ & new_n4844_;
  assign new_n4851_ = ~new_n4850_;
  assign new_n4852_ = new_n4851_ & new_n264_;
  assign new_n4853_ = ~new_n4852_;
  assign new_n4854_ = new_n3089_ & new_n369_;
  assign new_n4855_ = ~new_n4854_;
  assign new_n4856_ = new_n3103_ & new_n469_;
  assign new_n4857_ = ~new_n4856_;
  assign new_n4858_ = new_n4857_ & new_n4855_;
  assign new_n4859_ = new_n3041_ & new_n570_;
  assign new_n4860_ = ~new_n4859_;
  assign new_n4861_ = new_n3027_ & new_n669_;
  assign new_n4862_ = ~new_n4861_;
  assign new_n4863_ = new_n4862_ & new_n4860_;
  assign new_n4864_ = new_n4863_ & new_n4858_;
  assign new_n4865_ = ~new_n4864_;
  assign new_n4866_ = new_n4865_ & shift6;
  assign new_n4867_ = ~new_n4866_;
  assign new_n4868_ = new_n4867_ & new_n4853_;
  assign ores39 = ~new_n4868_;
  assign new_n4870_ = new_n3258_ & new_n669_;
  assign new_n4871_ = ~new_n4870_;
  assign new_n4872_ = new_n3244_ & new_n570_;
  assign new_n4873_ = ~new_n4872_;
  assign new_n4874_ = new_n4873_ & new_n4871_;
  assign new_n4875_ = new_n3182_ & new_n469_;
  assign new_n4876_ = ~new_n4875_;
  assign new_n4877_ = new_n3196_ & new_n369_;
  assign new_n4878_ = ~new_n4877_;
  assign new_n4879_ = new_n4878_ & new_n4876_;
  assign new_n4880_ = new_n4879_ & new_n4874_;
  assign new_n4881_ = ~new_n4880_;
  assign new_n4882_ = new_n4881_ & new_n264_;
  assign new_n4883_ = ~new_n4882_;
  assign new_n4884_ = new_n3215_ & new_n369_;
  assign new_n4885_ = ~new_n4884_;
  assign new_n4886_ = new_n3229_ & new_n469_;
  assign new_n4887_ = ~new_n4886_;
  assign new_n4888_ = new_n4887_ & new_n4885_;
  assign new_n4889_ = new_n3167_ & new_n570_;
  assign new_n4890_ = ~new_n4889_;
  assign new_n4891_ = new_n3153_ & new_n669_;
  assign new_n4892_ = ~new_n4891_;
  assign new_n4893_ = new_n4892_ & new_n4890_;
  assign new_n4894_ = new_n4893_ & new_n4888_;
  assign new_n4895_ = ~new_n4894_;
  assign new_n4896_ = new_n4895_ & shift6;
  assign new_n4897_ = ~new_n4896_;
  assign new_n4898_ = new_n4897_ & new_n4883_;
  assign ores40 = ~new_n4898_;
  assign new_n4900_ = new_n3384_ & new_n669_;
  assign new_n4901_ = ~new_n4900_;
  assign new_n4902_ = new_n3370_ & new_n570_;
  assign new_n4903_ = ~new_n4902_;
  assign new_n4904_ = new_n4903_ & new_n4901_;
  assign new_n4905_ = new_n3308_ & new_n469_;
  assign new_n4906_ = ~new_n4905_;
  assign new_n4907_ = new_n3322_ & new_n369_;
  assign new_n4908_ = ~new_n4907_;
  assign new_n4909_ = new_n4908_ & new_n4906_;
  assign new_n4910_ = new_n4909_ & new_n4904_;
  assign new_n4911_ = ~new_n4910_;
  assign new_n4912_ = new_n4911_ & new_n264_;
  assign new_n4913_ = ~new_n4912_;
  assign new_n4914_ = new_n3341_ & new_n369_;
  assign new_n4915_ = ~new_n4914_;
  assign new_n4916_ = new_n3355_ & new_n469_;
  assign new_n4917_ = ~new_n4916_;
  assign new_n4918_ = new_n4917_ & new_n4915_;
  assign new_n4919_ = new_n3293_ & new_n570_;
  assign new_n4920_ = ~new_n4919_;
  assign new_n4921_ = new_n3279_ & new_n669_;
  assign new_n4922_ = ~new_n4921_;
  assign new_n4923_ = new_n4922_ & new_n4920_;
  assign new_n4924_ = new_n4923_ & new_n4918_;
  assign new_n4925_ = ~new_n4924_;
  assign new_n4926_ = new_n4925_ & shift6;
  assign new_n4927_ = ~new_n4926_;
  assign new_n4928_ = new_n4927_ & new_n4913_;
  assign ores41 = ~new_n4928_;
  assign new_n4930_ = new_n3448_ & new_n369_;
  assign new_n4931_ = ~new_n4930_;
  assign new_n4932_ = new_n3434_ & new_n469_;
  assign new_n4933_ = ~new_n4932_;
  assign new_n4934_ = new_n4933_ & new_n4931_;
  assign new_n4935_ = new_n3496_ & new_n570_;
  assign new_n4936_ = ~new_n4935_;
  assign new_n4937_ = new_n3510_ & new_n669_;
  assign new_n4938_ = ~new_n4937_;
  assign new_n4939_ = new_n4938_ & new_n4936_;
  assign new_n4940_ = new_n4939_ & new_n4934_;
  assign new_n4941_ = ~new_n4940_;
  assign new_n4942_ = new_n4941_ & new_n264_;
  assign new_n4943_ = ~new_n4942_;
  assign new_n4944_ = new_n3467_ & new_n369_;
  assign new_n4945_ = ~new_n4944_;
  assign new_n4946_ = new_n3481_ & new_n469_;
  assign new_n4947_ = ~new_n4946_;
  assign new_n4948_ = new_n4947_ & new_n4945_;
  assign new_n4949_ = new_n3419_ & new_n570_;
  assign new_n4950_ = ~new_n4949_;
  assign new_n4951_ = new_n3405_ & new_n669_;
  assign new_n4952_ = ~new_n4951_;
  assign new_n4953_ = new_n4952_ & new_n4950_;
  assign new_n4954_ = new_n4953_ & new_n4948_;
  assign new_n4955_ = ~new_n4954_;
  assign new_n4956_ = new_n4955_ & shift6;
  assign new_n4957_ = ~new_n4956_;
  assign new_n4958_ = new_n4957_ & new_n4943_;
  assign ores42 = ~new_n4958_;
  assign new_n4960_ = new_n3574_ & new_n369_;
  assign new_n4961_ = ~new_n4960_;
  assign new_n4962_ = new_n3560_ & new_n469_;
  assign new_n4963_ = ~new_n4962_;
  assign new_n4964_ = new_n4963_ & new_n4961_;
  assign new_n4965_ = new_n3622_ & new_n570_;
  assign new_n4966_ = ~new_n4965_;
  assign new_n4967_ = new_n3636_ & new_n669_;
  assign new_n4968_ = ~new_n4967_;
  assign new_n4969_ = new_n4968_ & new_n4966_;
  assign new_n4970_ = new_n4969_ & new_n4964_;
  assign new_n4971_ = ~new_n4970_;
  assign new_n4972_ = new_n4971_ & new_n264_;
  assign new_n4973_ = ~new_n4972_;
  assign new_n4974_ = new_n3593_ & new_n369_;
  assign new_n4975_ = ~new_n4974_;
  assign new_n4976_ = new_n3607_ & new_n469_;
  assign new_n4977_ = ~new_n4976_;
  assign new_n4978_ = new_n4977_ & new_n4975_;
  assign new_n4979_ = new_n3545_ & new_n570_;
  assign new_n4980_ = ~new_n4979_;
  assign new_n4981_ = new_n3531_ & new_n669_;
  assign new_n4982_ = ~new_n4981_;
  assign new_n4983_ = new_n4982_ & new_n4980_;
  assign new_n4984_ = new_n4983_ & new_n4978_;
  assign new_n4985_ = ~new_n4984_;
  assign new_n4986_ = new_n4985_ & shift6;
  assign new_n4987_ = ~new_n4986_;
  assign new_n4988_ = new_n4987_ & new_n4973_;
  assign ores43 = ~new_n4988_;
  assign new_n4990_ = new_n3700_ & new_n369_;
  assign new_n4991_ = ~new_n4990_;
  assign new_n4992_ = new_n3686_ & new_n469_;
  assign new_n4993_ = ~new_n4992_;
  assign new_n4994_ = new_n4993_ & new_n4991_;
  assign new_n4995_ = new_n3748_ & new_n570_;
  assign new_n4996_ = ~new_n4995_;
  assign new_n4997_ = new_n3762_ & new_n669_;
  assign new_n4998_ = ~new_n4997_;
  assign new_n4999_ = new_n4998_ & new_n4996_;
  assign new_n5000_ = new_n4999_ & new_n4994_;
  assign new_n5001_ = ~new_n5000_;
  assign new_n5002_ = new_n5001_ & new_n264_;
  assign new_n5003_ = ~new_n5002_;
  assign new_n5004_ = new_n3719_ & new_n369_;
  assign new_n5005_ = ~new_n5004_;
  assign new_n5006_ = new_n3733_ & new_n469_;
  assign new_n5007_ = ~new_n5006_;
  assign new_n5008_ = new_n5007_ & new_n5005_;
  assign new_n5009_ = new_n3671_ & new_n570_;
  assign new_n5010_ = ~new_n5009_;
  assign new_n5011_ = new_n3657_ & new_n669_;
  assign new_n5012_ = ~new_n5011_;
  assign new_n5013_ = new_n5012_ & new_n5010_;
  assign new_n5014_ = new_n5013_ & new_n5008_;
  assign new_n5015_ = ~new_n5014_;
  assign new_n5016_ = new_n5015_ & shift6;
  assign new_n5017_ = ~new_n5016_;
  assign new_n5018_ = new_n5017_ & new_n5003_;
  assign ores44 = ~new_n5018_;
  assign new_n5020_ = new_n3826_ & new_n369_;
  assign new_n5021_ = ~new_n5020_;
  assign new_n5022_ = new_n3812_ & new_n469_;
  assign new_n5023_ = ~new_n5022_;
  assign new_n5024_ = new_n5023_ & new_n5021_;
  assign new_n5025_ = new_n3874_ & new_n570_;
  assign new_n5026_ = ~new_n5025_;
  assign new_n5027_ = new_n3888_ & new_n669_;
  assign new_n5028_ = ~new_n5027_;
  assign new_n5029_ = new_n5028_ & new_n5026_;
  assign new_n5030_ = new_n5029_ & new_n5024_;
  assign new_n5031_ = ~new_n5030_;
  assign new_n5032_ = new_n5031_ & new_n264_;
  assign new_n5033_ = ~new_n5032_;
  assign new_n5034_ = new_n3845_ & new_n369_;
  assign new_n5035_ = ~new_n5034_;
  assign new_n5036_ = new_n3859_ & new_n469_;
  assign new_n5037_ = ~new_n5036_;
  assign new_n5038_ = new_n5037_ & new_n5035_;
  assign new_n5039_ = new_n3797_ & new_n570_;
  assign new_n5040_ = ~new_n5039_;
  assign new_n5041_ = new_n3783_ & new_n669_;
  assign new_n5042_ = ~new_n5041_;
  assign new_n5043_ = new_n5042_ & new_n5040_;
  assign new_n5044_ = new_n5043_ & new_n5038_;
  assign new_n5045_ = ~new_n5044_;
  assign new_n5046_ = new_n5045_ & shift6;
  assign new_n5047_ = ~new_n5046_;
  assign new_n5048_ = new_n5047_ & new_n5033_;
  assign ores45 = ~new_n5048_;
  assign new_n5050_ = new_n3952_ & new_n369_;
  assign new_n5051_ = ~new_n5050_;
  assign new_n5052_ = new_n3938_ & new_n469_;
  assign new_n5053_ = ~new_n5052_;
  assign new_n5054_ = new_n5053_ & new_n5051_;
  assign new_n5055_ = new_n4000_ & new_n570_;
  assign new_n5056_ = ~new_n5055_;
  assign new_n5057_ = new_n4014_ & new_n669_;
  assign new_n5058_ = ~new_n5057_;
  assign new_n5059_ = new_n5058_ & new_n5056_;
  assign new_n5060_ = new_n5059_ & new_n5054_;
  assign new_n5061_ = ~new_n5060_;
  assign new_n5062_ = new_n5061_ & new_n264_;
  assign new_n5063_ = ~new_n5062_;
  assign new_n5064_ = new_n3971_ & new_n369_;
  assign new_n5065_ = ~new_n5064_;
  assign new_n5066_ = new_n3985_ & new_n469_;
  assign new_n5067_ = ~new_n5066_;
  assign new_n5068_ = new_n5067_ & new_n5065_;
  assign new_n5069_ = new_n3923_ & new_n570_;
  assign new_n5070_ = ~new_n5069_;
  assign new_n5071_ = new_n3909_ & new_n669_;
  assign new_n5072_ = ~new_n5071_;
  assign new_n5073_ = new_n5072_ & new_n5070_;
  assign new_n5074_ = new_n5073_ & new_n5068_;
  assign new_n5075_ = ~new_n5074_;
  assign new_n5076_ = new_n5075_ & shift6;
  assign new_n5077_ = ~new_n5076_;
  assign new_n5078_ = new_n5077_ & new_n5063_;
  assign ores46 = ~new_n5078_;
  assign new_n5080_ = new_n4078_ & new_n369_;
  assign new_n5081_ = ~new_n5080_;
  assign new_n5082_ = new_n4064_ & new_n469_;
  assign new_n5083_ = ~new_n5082_;
  assign new_n5084_ = new_n5083_ & new_n5081_;
  assign new_n5085_ = new_n4126_ & new_n570_;
  assign new_n5086_ = ~new_n5085_;
  assign new_n5087_ = new_n4140_ & new_n669_;
  assign new_n5088_ = ~new_n5087_;
  assign new_n5089_ = new_n5088_ & new_n5086_;
  assign new_n5090_ = new_n5089_ & new_n5084_;
  assign new_n5091_ = ~new_n5090_;
  assign new_n5092_ = new_n5091_ & new_n264_;
  assign new_n5093_ = ~new_n5092_;
  assign new_n5094_ = new_n4097_ & new_n369_;
  assign new_n5095_ = ~new_n5094_;
  assign new_n5096_ = new_n4111_ & new_n469_;
  assign new_n5097_ = ~new_n5096_;
  assign new_n5098_ = new_n5097_ & new_n5095_;
  assign new_n5099_ = new_n4049_ & new_n570_;
  assign new_n5100_ = ~new_n5099_;
  assign new_n5101_ = new_n4035_ & new_n669_;
  assign new_n5102_ = ~new_n5101_;
  assign new_n5103_ = new_n5102_ & new_n5100_;
  assign new_n5104_ = new_n5103_ & new_n5098_;
  assign new_n5105_ = ~new_n5104_;
  assign new_n5106_ = new_n5105_ & shift6;
  assign new_n5107_ = ~new_n5106_;
  assign new_n5108_ = new_n5107_ & new_n5093_;
  assign ores47 = ~new_n5108_;
  assign new_n5110_ = new_n568_ & new_n369_;
  assign new_n5111_ = ~new_n5110_;
  assign new_n5112_ = new_n772_ & new_n469_;
  assign new_n5113_ = ~new_n5112_;
  assign new_n5114_ = new_n5113_ & new_n5111_;
  assign new_n5115_ = new_n1065_ & new_n570_;
  assign new_n5116_ = ~new_n5115_;
  assign new_n5117_ = new_n870_ & new_n669_;
  assign new_n5118_ = ~new_n5117_;
  assign new_n5119_ = new_n5118_ & new_n5116_;
  assign new_n5120_ = new_n5119_ & new_n5114_;
  assign new_n5121_ = ~new_n5120_;
  assign new_n5122_ = new_n5121_ & new_n264_;
  assign new_n5123_ = ~new_n5122_;
  assign new_n5124_ = new_n469_ & new_n368_;
  assign new_n5125_ = ~new_n5124_;
  assign new_n5126_ = new_n669_ & new_n467_;
  assign new_n5127_ = ~new_n5126_;
  assign new_n5128_ = new_n5127_ & new_n5125_;
  assign new_n5129_ = new_n969_ & new_n369_;
  assign new_n5130_ = ~new_n5129_;
  assign new_n5131_ = new_n668_ & new_n570_;
  assign new_n5132_ = ~new_n5131_;
  assign new_n5133_ = new_n5132_ & new_n5130_;
  assign new_n5134_ = new_n5133_ & new_n5128_;
  assign new_n5135_ = ~new_n5134_;
  assign new_n5136_ = new_n5135_ & shift6;
  assign new_n5137_ = ~new_n5136_;
  assign new_n5138_ = new_n5137_ & new_n5123_;
  assign ores48 = ~new_n5138_;
  assign new_n5140_ = new_n1343_ & new_n369_;
  assign new_n5141_ = ~new_n5140_;
  assign new_n5142_ = new_n1618_ & new_n469_;
  assign new_n5143_ = ~new_n5142_;
  assign new_n5144_ = new_n5143_ & new_n5141_;
  assign new_n5145_ = new_n1706_ & new_n570_;
  assign new_n5146_ = ~new_n5145_;
  assign new_n5147_ = new_n1796_ & new_n669_;
  assign new_n5148_ = ~new_n5147_;
  assign new_n5149_ = new_n5148_ & new_n5146_;
  assign new_n5150_ = new_n5149_ & new_n5144_;
  assign new_n5151_ = ~new_n5150_;
  assign new_n5152_ = new_n5151_ & new_n264_;
  assign new_n5153_ = ~new_n5152_;
  assign new_n5154_ = new_n1528_ & new_n369_;
  assign new_n5155_ = ~new_n5154_;
  assign new_n5156_ = new_n1162_ & new_n469_;
  assign new_n5157_ = ~new_n5156_;
  assign new_n5158_ = new_n5157_ & new_n5155_;
  assign new_n5159_ = new_n1433_ & new_n570_;
  assign new_n5160_ = ~new_n5159_;
  assign new_n5161_ = new_n1252_ & new_n669_;
  assign new_n5162_ = ~new_n5161_;
  assign new_n5163_ = new_n5162_ & new_n5160_;
  assign new_n5164_ = new_n5163_ & new_n5158_;
  assign new_n5165_ = ~new_n5164_;
  assign new_n5166_ = new_n5165_ & shift6;
  assign new_n5167_ = ~new_n5166_;
  assign new_n5168_ = new_n5167_ & new_n5153_;
  assign ores49 = ~new_n5168_;
  assign new_n5170_ = new_n1906_ & new_n369_;
  assign new_n5171_ = ~new_n5170_;
  assign new_n5172_ = new_n2013_ & new_n469_;
  assign new_n5173_ = ~new_n5172_;
  assign new_n5174_ = new_n5173_ & new_n5171_;
  assign new_n5175_ = new_n2056_ & new_n570_;
  assign new_n5176_ = ~new_n5175_;
  assign new_n5177_ = new_n2090_ & new_n669_;
  assign new_n5178_ = ~new_n5177_;
  assign new_n5179_ = new_n5178_ & new_n5176_;
  assign new_n5180_ = new_n5179_ & new_n5174_;
  assign new_n5181_ = ~new_n5180_;
  assign new_n5182_ = new_n5181_ & new_n264_;
  assign new_n5183_ = ~new_n5182_;
  assign new_n5184_ = new_n1979_ & new_n369_;
  assign new_n5185_ = ~new_n5184_;
  assign new_n5186_ = new_n1837_ & new_n469_;
  assign new_n5187_ = ~new_n5186_;
  assign new_n5188_ = new_n5187_ & new_n5185_;
  assign new_n5189_ = new_n1940_ & new_n570_;
  assign new_n5190_ = ~new_n5189_;
  assign new_n5191_ = new_n1871_ & new_n669_;
  assign new_n5192_ = ~new_n5191_;
  assign new_n5193_ = new_n5192_ & new_n5190_;
  assign new_n5194_ = new_n5193_ & new_n5188_;
  assign new_n5195_ = ~new_n5194_;
  assign new_n5196_ = new_n5195_ & shift6;
  assign new_n5197_ = ~new_n5196_;
  assign new_n5198_ = new_n5197_ & new_n5183_;
  assign ores50 = ~new_n5198_;
  assign new_n5200_ = new_n2495_ & new_n570_;
  assign new_n5201_ = ~new_n5200_;
  assign new_n5202_ = new_n2628_ & new_n669_;
  assign new_n5203_ = ~new_n5202_;
  assign new_n5204_ = new_n5203_ & new_n5201_;
  assign new_n5205_ = new_n2296_ & new_n369_;
  assign new_n5206_ = ~new_n5205_;
  assign new_n5207_ = new_n2562_ & new_n469_;
  assign new_n5208_ = ~new_n5207_;
  assign new_n5209_ = new_n5208_ & new_n5206_;
  assign new_n5210_ = new_n5209_ & new_n5204_;
  assign new_n5211_ = ~new_n5210_;
  assign new_n5212_ = new_n5211_ & new_n264_;
  assign new_n5213_ = ~new_n5212_;
  assign new_n5214_ = new_n2433_ & new_n369_;
  assign new_n5215_ = ~new_n5214_;
  assign new_n5216_ = new_n2163_ & new_n570_;
  assign new_n5217_ = ~new_n5216_;
  assign new_n5218_ = new_n5217_ & new_n5215_;
  assign new_n5219_ = new_n2362_ & new_n469_;
  assign new_n5220_ = ~new_n5219_;
  assign new_n5221_ = new_n2229_ & new_n669_;
  assign new_n5222_ = ~new_n5221_;
  assign new_n5223_ = new_n5222_ & new_n5220_;
  assign new_n5224_ = new_n5223_ & new_n5218_;
  assign new_n5225_ = ~new_n5224_;
  assign new_n5226_ = new_n5225_ & shift6;
  assign new_n5227_ = ~new_n5226_;
  assign new_n5228_ = new_n5227_ & new_n5213_;
  assign ores51 = ~new_n5228_;
  assign new_n5230_ = new_n2711_ & new_n570_;
  assign new_n5231_ = ~new_n5230_;
  assign new_n5232_ = new_n2678_ & new_n369_;
  assign new_n5233_ = ~new_n5232_;
  assign new_n5234_ = new_n5233_ & new_n5231_;
  assign new_n5235_ = new_n2740_ & new_n669_;
  assign new_n5236_ = ~new_n5235_;
  assign new_n5237_ = new_n2754_ & new_n469_;
  assign new_n5238_ = ~new_n5237_;
  assign new_n5239_ = new_n5238_ & new_n5236_;
  assign new_n5240_ = new_n5239_ & new_n5234_;
  assign new_n5241_ = ~new_n5240_;
  assign new_n5242_ = new_n5241_ & new_n264_;
  assign new_n5243_ = ~new_n5242_;
  assign new_n5244_ = new_n2649_ & new_n469_;
  assign new_n5245_ = ~new_n5244_;
  assign new_n5246_ = new_n2663_ & new_n669_;
  assign new_n5247_ = ~new_n5246_;
  assign new_n5248_ = new_n5247_ & new_n5245_;
  assign new_n5249_ = new_n2692_ & new_n570_;
  assign new_n5250_ = ~new_n5249_;
  assign new_n5251_ = new_n2725_ & new_n369_;
  assign new_n5252_ = ~new_n5251_;
  assign new_n5253_ = new_n5252_ & new_n5250_;
  assign new_n5254_ = new_n5253_ & new_n5248_;
  assign new_n5255_ = ~new_n5254_;
  assign new_n5256_ = new_n5255_ & shift6;
  assign new_n5257_ = ~new_n5256_;
  assign new_n5258_ = new_n5257_ & new_n5243_;
  assign ores52 = ~new_n5258_;
  assign new_n5260_ = new_n2837_ & new_n570_;
  assign new_n5261_ = ~new_n5260_;
  assign new_n5262_ = new_n2804_ & new_n369_;
  assign new_n5263_ = ~new_n5262_;
  assign new_n5264_ = new_n5263_ & new_n5261_;
  assign new_n5265_ = new_n2866_ & new_n669_;
  assign new_n5266_ = ~new_n5265_;
  assign new_n5267_ = new_n2880_ & new_n469_;
  assign new_n5268_ = ~new_n5267_;
  assign new_n5269_ = new_n5268_ & new_n5266_;
  assign new_n5270_ = new_n5269_ & new_n5264_;
  assign new_n5271_ = ~new_n5270_;
  assign new_n5272_ = new_n5271_ & new_n264_;
  assign new_n5273_ = ~new_n5272_;
  assign new_n5274_ = new_n2775_ & new_n469_;
  assign new_n5275_ = ~new_n5274_;
  assign new_n5276_ = new_n2789_ & new_n669_;
  assign new_n5277_ = ~new_n5276_;
  assign new_n5278_ = new_n5277_ & new_n5275_;
  assign new_n5279_ = new_n2818_ & new_n570_;
  assign new_n5280_ = ~new_n5279_;
  assign new_n5281_ = new_n2851_ & new_n369_;
  assign new_n5282_ = ~new_n5281_;
  assign new_n5283_ = new_n5282_ & new_n5280_;
  assign new_n5284_ = new_n5283_ & new_n5278_;
  assign new_n5285_ = ~new_n5284_;
  assign new_n5286_ = new_n5285_ & shift6;
  assign new_n5287_ = ~new_n5286_;
  assign new_n5288_ = new_n5287_ & new_n5273_;
  assign ores53 = ~new_n5288_;
  assign new_n5290_ = new_n2963_ & new_n570_;
  assign new_n5291_ = ~new_n5290_;
  assign new_n5292_ = new_n2930_ & new_n369_;
  assign new_n5293_ = ~new_n5292_;
  assign new_n5294_ = new_n5293_ & new_n5291_;
  assign new_n5295_ = new_n2992_ & new_n669_;
  assign new_n5296_ = ~new_n5295_;
  assign new_n5297_ = new_n3006_ & new_n469_;
  assign new_n5298_ = ~new_n5297_;
  assign new_n5299_ = new_n5298_ & new_n5296_;
  assign new_n5300_ = new_n5299_ & new_n5294_;
  assign new_n5301_ = ~new_n5300_;
  assign new_n5302_ = new_n5301_ & new_n264_;
  assign new_n5303_ = ~new_n5302_;
  assign new_n5304_ = new_n2901_ & new_n469_;
  assign new_n5305_ = ~new_n5304_;
  assign new_n5306_ = new_n2915_ & new_n669_;
  assign new_n5307_ = ~new_n5306_;
  assign new_n5308_ = new_n5307_ & new_n5305_;
  assign new_n5309_ = new_n2944_ & new_n570_;
  assign new_n5310_ = ~new_n5309_;
  assign new_n5311_ = new_n2977_ & new_n369_;
  assign new_n5312_ = ~new_n5311_;
  assign new_n5313_ = new_n5312_ & new_n5310_;
  assign new_n5314_ = new_n5313_ & new_n5308_;
  assign new_n5315_ = ~new_n5314_;
  assign new_n5316_ = new_n5315_ & shift6;
  assign new_n5317_ = ~new_n5316_;
  assign new_n5318_ = new_n5317_ & new_n5303_;
  assign ores54 = ~new_n5318_;
  assign new_n5320_ = new_n3089_ & new_n570_;
  assign new_n5321_ = ~new_n5320_;
  assign new_n5322_ = new_n3132_ & new_n469_;
  assign new_n5323_ = ~new_n5322_;
  assign new_n5324_ = new_n5323_ & new_n5321_;
  assign new_n5325_ = new_n3056_ & new_n369_;
  assign new_n5326_ = ~new_n5325_;
  assign new_n5327_ = new_n3118_ & new_n669_;
  assign new_n5328_ = ~new_n5327_;
  assign new_n5329_ = new_n5328_ & new_n5326_;
  assign new_n5330_ = new_n5329_ & new_n5324_;
  assign new_n5331_ = ~new_n5330_;
  assign new_n5332_ = new_n5331_ & new_n264_;
  assign new_n5333_ = ~new_n5332_;
  assign new_n5334_ = new_n3103_ & new_n369_;
  assign new_n5335_ = ~new_n5334_;
  assign new_n5336_ = new_n3027_ & new_n469_;
  assign new_n5337_ = ~new_n5336_;
  assign new_n5338_ = new_n5337_ & new_n5335_;
  assign new_n5339_ = new_n3070_ & new_n570_;
  assign new_n5340_ = ~new_n5339_;
  assign new_n5341_ = new_n3041_ & new_n669_;
  assign new_n5342_ = ~new_n5341_;
  assign new_n5343_ = new_n5342_ & new_n5340_;
  assign new_n5344_ = new_n5343_ & new_n5338_;
  assign new_n5345_ = ~new_n5344_;
  assign new_n5346_ = new_n5345_ & shift6;
  assign new_n5347_ = ~new_n5346_;
  assign new_n5348_ = new_n5347_ & new_n5333_;
  assign ores55 = ~new_n5348_;
  assign new_n5350_ = new_n3215_ & new_n570_;
  assign new_n5351_ = ~new_n5350_;
  assign new_n5352_ = new_n3258_ & new_n469_;
  assign new_n5353_ = ~new_n5352_;
  assign new_n5354_ = new_n5353_ & new_n5351_;
  assign new_n5355_ = new_n3182_ & new_n369_;
  assign new_n5356_ = ~new_n5355_;
  assign new_n5357_ = new_n3244_ & new_n669_;
  assign new_n5358_ = ~new_n5357_;
  assign new_n5359_ = new_n5358_ & new_n5356_;
  assign new_n5360_ = new_n5359_ & new_n5354_;
  assign new_n5361_ = ~new_n5360_;
  assign new_n5362_ = new_n5361_ & new_n264_;
  assign new_n5363_ = ~new_n5362_;
  assign new_n5364_ = new_n3229_ & new_n369_;
  assign new_n5365_ = ~new_n5364_;
  assign new_n5366_ = new_n3153_ & new_n469_;
  assign new_n5367_ = ~new_n5366_;
  assign new_n5368_ = new_n5367_ & new_n5365_;
  assign new_n5369_ = new_n3196_ & new_n570_;
  assign new_n5370_ = ~new_n5369_;
  assign new_n5371_ = new_n3167_ & new_n669_;
  assign new_n5372_ = ~new_n5371_;
  assign new_n5373_ = new_n5372_ & new_n5370_;
  assign new_n5374_ = new_n5373_ & new_n5368_;
  assign new_n5375_ = ~new_n5374_;
  assign new_n5376_ = new_n5375_ & shift6;
  assign new_n5377_ = ~new_n5376_;
  assign new_n5378_ = new_n5377_ & new_n5363_;
  assign ores56 = ~new_n5378_;
  assign new_n5380_ = new_n3341_ & new_n570_;
  assign new_n5381_ = ~new_n5380_;
  assign new_n5382_ = new_n3384_ & new_n469_;
  assign new_n5383_ = ~new_n5382_;
  assign new_n5384_ = new_n5383_ & new_n5381_;
  assign new_n5385_ = new_n3308_ & new_n369_;
  assign new_n5386_ = ~new_n5385_;
  assign new_n5387_ = new_n3370_ & new_n669_;
  assign new_n5388_ = ~new_n5387_;
  assign new_n5389_ = new_n5388_ & new_n5386_;
  assign new_n5390_ = new_n5389_ & new_n5384_;
  assign new_n5391_ = ~new_n5390_;
  assign new_n5392_ = new_n5391_ & new_n264_;
  assign new_n5393_ = ~new_n5392_;
  assign new_n5394_ = new_n3355_ & new_n369_;
  assign new_n5395_ = ~new_n5394_;
  assign new_n5396_ = new_n3279_ & new_n469_;
  assign new_n5397_ = ~new_n5396_;
  assign new_n5398_ = new_n5397_ & new_n5395_;
  assign new_n5399_ = new_n3322_ & new_n570_;
  assign new_n5400_ = ~new_n5399_;
  assign new_n5401_ = new_n3293_ & new_n669_;
  assign new_n5402_ = ~new_n5401_;
  assign new_n5403_ = new_n5402_ & new_n5400_;
  assign new_n5404_ = new_n5403_ & new_n5398_;
  assign new_n5405_ = ~new_n5404_;
  assign new_n5406_ = new_n5405_ & shift6;
  assign new_n5407_ = ~new_n5406_;
  assign new_n5408_ = new_n5407_ & new_n5393_;
  assign ores57 = ~new_n5408_;
  assign new_n5410_ = new_n3467_ & new_n570_;
  assign new_n5411_ = ~new_n5410_;
  assign new_n5412_ = new_n3434_ & new_n369_;
  assign new_n5413_ = ~new_n5412_;
  assign new_n5414_ = new_n5413_ & new_n5411_;
  assign new_n5415_ = new_n3496_ & new_n669_;
  assign new_n5416_ = ~new_n5415_;
  assign new_n5417_ = new_n3510_ & new_n469_;
  assign new_n5418_ = ~new_n5417_;
  assign new_n5419_ = new_n5418_ & new_n5416_;
  assign new_n5420_ = new_n5419_ & new_n5414_;
  assign new_n5421_ = ~new_n5420_;
  assign new_n5422_ = new_n5421_ & new_n264_;
  assign new_n5423_ = ~new_n5422_;
  assign new_n5424_ = new_n3481_ & new_n369_;
  assign new_n5425_ = ~new_n5424_;
  assign new_n5426_ = new_n3405_ & new_n469_;
  assign new_n5427_ = ~new_n5426_;
  assign new_n5428_ = new_n5427_ & new_n5425_;
  assign new_n5429_ = new_n3448_ & new_n570_;
  assign new_n5430_ = ~new_n5429_;
  assign new_n5431_ = new_n3419_ & new_n669_;
  assign new_n5432_ = ~new_n5431_;
  assign new_n5433_ = new_n5432_ & new_n5430_;
  assign new_n5434_ = new_n5433_ & new_n5428_;
  assign new_n5435_ = ~new_n5434_;
  assign new_n5436_ = new_n5435_ & shift6;
  assign new_n5437_ = ~new_n5436_;
  assign new_n5438_ = new_n5437_ & new_n5423_;
  assign ores58 = ~new_n5438_;
  assign new_n5440_ = new_n3593_ & new_n570_;
  assign new_n5441_ = ~new_n5440_;
  assign new_n5442_ = new_n3560_ & new_n369_;
  assign new_n5443_ = ~new_n5442_;
  assign new_n5444_ = new_n5443_ & new_n5441_;
  assign new_n5445_ = new_n3622_ & new_n669_;
  assign new_n5446_ = ~new_n5445_;
  assign new_n5447_ = new_n3636_ & new_n469_;
  assign new_n5448_ = ~new_n5447_;
  assign new_n5449_ = new_n5448_ & new_n5446_;
  assign new_n5450_ = new_n5449_ & new_n5444_;
  assign new_n5451_ = ~new_n5450_;
  assign new_n5452_ = new_n5451_ & new_n264_;
  assign new_n5453_ = ~new_n5452_;
  assign new_n5454_ = new_n3607_ & new_n369_;
  assign new_n5455_ = ~new_n5454_;
  assign new_n5456_ = new_n3531_ & new_n469_;
  assign new_n5457_ = ~new_n5456_;
  assign new_n5458_ = new_n5457_ & new_n5455_;
  assign new_n5459_ = new_n3574_ & new_n570_;
  assign new_n5460_ = ~new_n5459_;
  assign new_n5461_ = new_n3545_ & new_n669_;
  assign new_n5462_ = ~new_n5461_;
  assign new_n5463_ = new_n5462_ & new_n5460_;
  assign new_n5464_ = new_n5463_ & new_n5458_;
  assign new_n5465_ = ~new_n5464_;
  assign new_n5466_ = new_n5465_ & shift6;
  assign new_n5467_ = ~new_n5466_;
  assign new_n5468_ = new_n5467_ & new_n5453_;
  assign ores59 = ~new_n5468_;
  assign new_n5470_ = new_n3719_ & new_n570_;
  assign new_n5471_ = ~new_n5470_;
  assign new_n5472_ = new_n3686_ & new_n369_;
  assign new_n5473_ = ~new_n5472_;
  assign new_n5474_ = new_n5473_ & new_n5471_;
  assign new_n5475_ = new_n3748_ & new_n669_;
  assign new_n5476_ = ~new_n5475_;
  assign new_n5477_ = new_n3762_ & new_n469_;
  assign new_n5478_ = ~new_n5477_;
  assign new_n5479_ = new_n5478_ & new_n5476_;
  assign new_n5480_ = new_n5479_ & new_n5474_;
  assign new_n5481_ = ~new_n5480_;
  assign new_n5482_ = new_n5481_ & new_n264_;
  assign new_n5483_ = ~new_n5482_;
  assign new_n5484_ = new_n3733_ & new_n369_;
  assign new_n5485_ = ~new_n5484_;
  assign new_n5486_ = new_n3657_ & new_n469_;
  assign new_n5487_ = ~new_n5486_;
  assign new_n5488_ = new_n5487_ & new_n5485_;
  assign new_n5489_ = new_n3700_ & new_n570_;
  assign new_n5490_ = ~new_n5489_;
  assign new_n5491_ = new_n3671_ & new_n669_;
  assign new_n5492_ = ~new_n5491_;
  assign new_n5493_ = new_n5492_ & new_n5490_;
  assign new_n5494_ = new_n5493_ & new_n5488_;
  assign new_n5495_ = ~new_n5494_;
  assign new_n5496_ = new_n5495_ & shift6;
  assign new_n5497_ = ~new_n5496_;
  assign new_n5498_ = new_n5497_ & new_n5483_;
  assign ores60 = ~new_n5498_;
  assign new_n5500_ = new_n3845_ & new_n570_;
  assign new_n5501_ = ~new_n5500_;
  assign new_n5502_ = new_n3812_ & new_n369_;
  assign new_n5503_ = ~new_n5502_;
  assign new_n5504_ = new_n5503_ & new_n5501_;
  assign new_n5505_ = new_n3874_ & new_n669_;
  assign new_n5506_ = ~new_n5505_;
  assign new_n5507_ = new_n3888_ & new_n469_;
  assign new_n5508_ = ~new_n5507_;
  assign new_n5509_ = new_n5508_ & new_n5506_;
  assign new_n5510_ = new_n5509_ & new_n5504_;
  assign new_n5511_ = ~new_n5510_;
  assign new_n5512_ = new_n5511_ & new_n264_;
  assign new_n5513_ = ~new_n5512_;
  assign new_n5514_ = new_n3859_ & new_n369_;
  assign new_n5515_ = ~new_n5514_;
  assign new_n5516_ = new_n3783_ & new_n469_;
  assign new_n5517_ = ~new_n5516_;
  assign new_n5518_ = new_n5517_ & new_n5515_;
  assign new_n5519_ = new_n3826_ & new_n570_;
  assign new_n5520_ = ~new_n5519_;
  assign new_n5521_ = new_n3797_ & new_n669_;
  assign new_n5522_ = ~new_n5521_;
  assign new_n5523_ = new_n5522_ & new_n5520_;
  assign new_n5524_ = new_n5523_ & new_n5518_;
  assign new_n5525_ = ~new_n5524_;
  assign new_n5526_ = new_n5525_ & shift6;
  assign new_n5527_ = ~new_n5526_;
  assign new_n5528_ = new_n5527_ & new_n5513_;
  assign ores61 = ~new_n5528_;
  assign new_n5530_ = new_n3971_ & new_n570_;
  assign new_n5531_ = ~new_n5530_;
  assign new_n5532_ = new_n3938_ & new_n369_;
  assign new_n5533_ = ~new_n5532_;
  assign new_n5534_ = new_n5533_ & new_n5531_;
  assign new_n5535_ = new_n4000_ & new_n669_;
  assign new_n5536_ = ~new_n5535_;
  assign new_n5537_ = new_n4014_ & new_n469_;
  assign new_n5538_ = ~new_n5537_;
  assign new_n5539_ = new_n5538_ & new_n5536_;
  assign new_n5540_ = new_n5539_ & new_n5534_;
  assign new_n5541_ = ~new_n5540_;
  assign new_n5542_ = new_n5541_ & new_n264_;
  assign new_n5543_ = ~new_n5542_;
  assign new_n5544_ = new_n3985_ & new_n369_;
  assign new_n5545_ = ~new_n5544_;
  assign new_n5546_ = new_n3909_ & new_n469_;
  assign new_n5547_ = ~new_n5546_;
  assign new_n5548_ = new_n5547_ & new_n5545_;
  assign new_n5549_ = new_n3952_ & new_n570_;
  assign new_n5550_ = ~new_n5549_;
  assign new_n5551_ = new_n3923_ & new_n669_;
  assign new_n5552_ = ~new_n5551_;
  assign new_n5553_ = new_n5552_ & new_n5550_;
  assign new_n5554_ = new_n5553_ & new_n5548_;
  assign new_n5555_ = ~new_n5554_;
  assign new_n5556_ = new_n5555_ & shift6;
  assign new_n5557_ = ~new_n5556_;
  assign new_n5558_ = new_n5557_ & new_n5543_;
  assign ores62 = ~new_n5558_;
  assign new_n5560_ = new_n4097_ & new_n570_;
  assign new_n5561_ = ~new_n5560_;
  assign new_n5562_ = new_n4064_ & new_n369_;
  assign new_n5563_ = ~new_n5562_;
  assign new_n5564_ = new_n5563_ & new_n5561_;
  assign new_n5565_ = new_n4126_ & new_n669_;
  assign new_n5566_ = ~new_n5565_;
  assign new_n5567_ = new_n4140_ & new_n469_;
  assign new_n5568_ = ~new_n5567_;
  assign new_n5569_ = new_n5568_ & new_n5566_;
  assign new_n5570_ = new_n5569_ & new_n5564_;
  assign new_n5571_ = ~new_n5570_;
  assign new_n5572_ = new_n5571_ & new_n264_;
  assign new_n5573_ = ~new_n5572_;
  assign new_n5574_ = new_n4111_ & new_n369_;
  assign new_n5575_ = ~new_n5574_;
  assign new_n5576_ = new_n4035_ & new_n469_;
  assign new_n5577_ = ~new_n5576_;
  assign new_n5578_ = new_n5577_ & new_n5575_;
  assign new_n5579_ = new_n4078_ & new_n570_;
  assign new_n5580_ = ~new_n5579_;
  assign new_n5581_ = new_n4049_ & new_n669_;
  assign new_n5582_ = ~new_n5581_;
  assign new_n5583_ = new_n5582_ & new_n5580_;
  assign new_n5584_ = new_n5583_ & new_n5578_;
  assign new_n5585_ = ~new_n5584_;
  assign new_n5586_ = new_n5585_ & shift6;
  assign new_n5587_ = ~new_n5586_;
  assign new_n5588_ = new_n5587_ & new_n5573_;
  assign ores63 = ~new_n5588_;
  assign new_n5590_ = new_n1070_ & new_n264_;
  assign new_n5591_ = ~new_n5590_;
  assign new_n5592_ = new_n674_ & shift6;
  assign new_n5593_ = ~new_n5592_;
  assign new_n5594_ = new_n5593_ & new_n5591_;
  assign ores64 = ~new_n5594_;
  assign new_n5596_ = new_n1801_ & new_n264_;
  assign new_n5597_ = ~new_n5596_;
  assign new_n5598_ = new_n1438_ & shift6;
  assign new_n5599_ = ~new_n5598_;
  assign new_n5600_ = new_n5599_ & new_n5597_;
  assign ores65 = ~new_n5600_;
  assign new_n5602_ = new_n2095_ & new_n264_;
  assign new_n5603_ = ~new_n5602_;
  assign new_n5604_ = new_n1945_ & shift6;
  assign new_n5605_ = ~new_n5604_;
  assign new_n5606_ = new_n5605_ & new_n5603_;
  assign ores66 = ~new_n5606_;
  assign new_n5608_ = new_n2633_ & new_n264_;
  assign new_n5609_ = ~new_n5608_;
  assign new_n5610_ = new_n2367_ & shift6;
  assign new_n5611_ = ~new_n5610_;
  assign new_n5612_ = new_n5611_ & new_n5609_;
  assign ores67 = ~new_n5612_;
  assign new_n5614_ = new_n2759_ & new_n264_;
  assign new_n5615_ = ~new_n5614_;
  assign new_n5616_ = new_n2697_ & shift6;
  assign new_n5617_ = ~new_n5616_;
  assign new_n5618_ = new_n5617_ & new_n5615_;
  assign ores68 = ~new_n5618_;
  assign new_n5620_ = new_n2885_ & new_n264_;
  assign new_n5621_ = ~new_n5620_;
  assign new_n5622_ = new_n2823_ & shift6;
  assign new_n5623_ = ~new_n5622_;
  assign new_n5624_ = new_n5623_ & new_n5621_;
  assign ores69 = ~new_n5624_;
  assign new_n5626_ = new_n3011_ & new_n264_;
  assign new_n5627_ = ~new_n5626_;
  assign new_n5628_ = new_n2949_ & shift6;
  assign new_n5629_ = ~new_n5628_;
  assign new_n5630_ = new_n5629_ & new_n5627_;
  assign ores70 = ~new_n5630_;
  assign new_n5632_ = new_n3137_ & new_n264_;
  assign new_n5633_ = ~new_n5632_;
  assign new_n5634_ = new_n3075_ & shift6;
  assign new_n5635_ = ~new_n5634_;
  assign new_n5636_ = new_n5635_ & new_n5633_;
  assign ores71 = ~new_n5636_;
  assign new_n5638_ = new_n3263_ & new_n264_;
  assign new_n5639_ = ~new_n5638_;
  assign new_n5640_ = new_n3201_ & shift6;
  assign new_n5641_ = ~new_n5640_;
  assign new_n5642_ = new_n5641_ & new_n5639_;
  assign ores72 = ~new_n5642_;
  assign new_n5644_ = new_n3389_ & new_n264_;
  assign new_n5645_ = ~new_n5644_;
  assign new_n5646_ = new_n3327_ & shift6;
  assign new_n5647_ = ~new_n5646_;
  assign new_n5648_ = new_n5647_ & new_n5645_;
  assign ores73 = ~new_n5648_;
  assign new_n5650_ = new_n3515_ & new_n264_;
  assign new_n5651_ = ~new_n5650_;
  assign new_n5652_ = new_n3453_ & shift6;
  assign new_n5653_ = ~new_n5652_;
  assign new_n5654_ = new_n5653_ & new_n5651_;
  assign ores74 = ~new_n5654_;
  assign new_n5656_ = new_n3641_ & new_n264_;
  assign new_n5657_ = ~new_n5656_;
  assign new_n5658_ = new_n3579_ & shift6;
  assign new_n5659_ = ~new_n5658_;
  assign new_n5660_ = new_n5659_ & new_n5657_;
  assign ores75 = ~new_n5660_;
  assign new_n5662_ = new_n3767_ & new_n264_;
  assign new_n5663_ = ~new_n5662_;
  assign new_n5664_ = new_n3705_ & shift6;
  assign new_n5665_ = ~new_n5664_;
  assign new_n5666_ = new_n5665_ & new_n5663_;
  assign ores76 = ~new_n5666_;
  assign new_n5668_ = new_n3893_ & new_n264_;
  assign new_n5669_ = ~new_n5668_;
  assign new_n5670_ = new_n3831_ & shift6;
  assign new_n5671_ = ~new_n5670_;
  assign new_n5672_ = new_n5671_ & new_n5669_;
  assign ores77 = ~new_n5672_;
  assign new_n5674_ = new_n4019_ & new_n264_;
  assign new_n5675_ = ~new_n5674_;
  assign new_n5676_ = new_n3957_ & shift6;
  assign new_n5677_ = ~new_n5676_;
  assign new_n5678_ = new_n5677_ & new_n5675_;
  assign ores78 = ~new_n5678_;
  assign new_n5680_ = new_n4145_ & new_n264_;
  assign new_n5681_ = ~new_n5680_;
  assign new_n5682_ = new_n4083_ & shift6;
  assign new_n5683_ = ~new_n5682_;
  assign new_n5684_ = new_n5683_ & new_n5681_;
  assign ores79 = ~new_n5684_;
  assign new_n5686_ = new_n4175_ & new_n264_;
  assign new_n5687_ = ~new_n5686_;
  assign new_n5688_ = new_n4161_ & shift6;
  assign new_n5689_ = ~new_n5688_;
  assign new_n5690_ = new_n5689_ & new_n5687_;
  assign ores80 = ~new_n5690_;
  assign new_n5692_ = new_n4205_ & new_n264_;
  assign new_n5693_ = ~new_n5692_;
  assign new_n5694_ = new_n4191_ & shift6;
  assign new_n5695_ = ~new_n5694_;
  assign new_n5696_ = new_n5695_ & new_n5693_;
  assign ores81 = ~new_n5696_;
  assign new_n5698_ = new_n4235_ & new_n264_;
  assign new_n5699_ = ~new_n5698_;
  assign new_n5700_ = new_n4221_ & shift6;
  assign new_n5701_ = ~new_n5700_;
  assign new_n5702_ = new_n5701_ & new_n5699_;
  assign ores82 = ~new_n5702_;
  assign new_n5704_ = new_n4265_ & new_n264_;
  assign new_n5705_ = ~new_n5704_;
  assign new_n5706_ = new_n4251_ & shift6;
  assign new_n5707_ = ~new_n5706_;
  assign new_n5708_ = new_n5707_ & new_n5705_;
  assign ores83 = ~new_n5708_;
  assign new_n5710_ = new_n4295_ & new_n264_;
  assign new_n5711_ = ~new_n5710_;
  assign new_n5712_ = new_n4281_ & shift6;
  assign new_n5713_ = ~new_n5712_;
  assign new_n5714_ = new_n5713_ & new_n5711_;
  assign ores84 = ~new_n5714_;
  assign new_n5716_ = new_n4325_ & new_n264_;
  assign new_n5717_ = ~new_n5716_;
  assign new_n5718_ = new_n4311_ & shift6;
  assign new_n5719_ = ~new_n5718_;
  assign new_n5720_ = new_n5719_ & new_n5717_;
  assign ores85 = ~new_n5720_;
  assign new_n5722_ = new_n4355_ & new_n264_;
  assign new_n5723_ = ~new_n5722_;
  assign new_n5724_ = new_n4341_ & shift6;
  assign new_n5725_ = ~new_n5724_;
  assign new_n5726_ = new_n5725_ & new_n5723_;
  assign ores86 = ~new_n5726_;
  assign new_n5728_ = new_n4385_ & new_n264_;
  assign new_n5729_ = ~new_n5728_;
  assign new_n5730_ = new_n4371_ & shift6;
  assign new_n5731_ = ~new_n5730_;
  assign new_n5732_ = new_n5731_ & new_n5729_;
  assign ores87 = ~new_n5732_;
  assign new_n5734_ = new_n4415_ & new_n264_;
  assign new_n5735_ = ~new_n5734_;
  assign new_n5736_ = new_n4401_ & shift6;
  assign new_n5737_ = ~new_n5736_;
  assign new_n5738_ = new_n5737_ & new_n5735_;
  assign ores88 = ~new_n5738_;
  assign new_n5740_ = new_n4445_ & new_n264_;
  assign new_n5741_ = ~new_n5740_;
  assign new_n5742_ = new_n4431_ & shift6;
  assign new_n5743_ = ~new_n5742_;
  assign new_n5744_ = new_n5743_ & new_n5741_;
  assign ores89 = ~new_n5744_;
  assign new_n5746_ = new_n4475_ & new_n264_;
  assign new_n5747_ = ~new_n5746_;
  assign new_n5748_ = new_n4461_ & shift6;
  assign new_n5749_ = ~new_n5748_;
  assign new_n5750_ = new_n5749_ & new_n5747_;
  assign ores90 = ~new_n5750_;
  assign new_n5752_ = new_n4505_ & new_n264_;
  assign new_n5753_ = ~new_n5752_;
  assign new_n5754_ = new_n4491_ & shift6;
  assign new_n5755_ = ~new_n5754_;
  assign new_n5756_ = new_n5755_ & new_n5753_;
  assign ores91 = ~new_n5756_;
  assign new_n5758_ = new_n4535_ & new_n264_;
  assign new_n5759_ = ~new_n5758_;
  assign new_n5760_ = new_n4521_ & shift6;
  assign new_n5761_ = ~new_n5760_;
  assign new_n5762_ = new_n5761_ & new_n5759_;
  assign ores92 = ~new_n5762_;
  assign new_n5764_ = new_n4565_ & new_n264_;
  assign new_n5765_ = ~new_n5764_;
  assign new_n5766_ = new_n4551_ & shift6;
  assign new_n5767_ = ~new_n5766_;
  assign new_n5768_ = new_n5767_ & new_n5765_;
  assign ores93 = ~new_n5768_;
  assign new_n5770_ = new_n4595_ & new_n264_;
  assign new_n5771_ = ~new_n5770_;
  assign new_n5772_ = new_n4581_ & shift6;
  assign new_n5773_ = ~new_n5772_;
  assign new_n5774_ = new_n5773_ & new_n5771_;
  assign ores94 = ~new_n5774_;
  assign new_n5776_ = new_n4625_ & new_n264_;
  assign new_n5777_ = ~new_n5776_;
  assign new_n5778_ = new_n4611_ & shift6;
  assign new_n5779_ = ~new_n5778_;
  assign new_n5780_ = new_n5779_ & new_n5777_;
  assign ores95 = ~new_n5780_;
  assign new_n5782_ = new_n4655_ & new_n264_;
  assign new_n5783_ = ~new_n5782_;
  assign new_n5784_ = new_n4641_ & shift6;
  assign new_n5785_ = ~new_n5784_;
  assign new_n5786_ = new_n5785_ & new_n5783_;
  assign ores96 = ~new_n5786_;
  assign new_n5788_ = new_n4685_ & new_n264_;
  assign new_n5789_ = ~new_n5788_;
  assign new_n5790_ = new_n4671_ & shift6;
  assign new_n5791_ = ~new_n5790_;
  assign new_n5792_ = new_n5791_ & new_n5789_;
  assign ores97 = ~new_n5792_;
  assign new_n5794_ = new_n4715_ & new_n264_;
  assign new_n5795_ = ~new_n5794_;
  assign new_n5796_ = new_n4701_ & shift6;
  assign new_n5797_ = ~new_n5796_;
  assign new_n5798_ = new_n5797_ & new_n5795_;
  assign ores98 = ~new_n5798_;
  assign new_n5800_ = new_n4745_ & new_n264_;
  assign new_n5801_ = ~new_n5800_;
  assign new_n5802_ = new_n4731_ & shift6;
  assign new_n5803_ = ~new_n5802_;
  assign new_n5804_ = new_n5803_ & new_n5801_;
  assign ores99 = ~new_n5804_;
  assign new_n5806_ = new_n4775_ & new_n264_;
  assign new_n5807_ = ~new_n5806_;
  assign new_n5808_ = new_n4761_ & shift6;
  assign new_n5809_ = ~new_n5808_;
  assign new_n5810_ = new_n5809_ & new_n5807_;
  assign ores100 = ~new_n5810_;
  assign new_n5812_ = new_n4805_ & new_n264_;
  assign new_n5813_ = ~new_n5812_;
  assign new_n5814_ = new_n4791_ & shift6;
  assign new_n5815_ = ~new_n5814_;
  assign new_n5816_ = new_n5815_ & new_n5813_;
  assign ores101 = ~new_n5816_;
  assign new_n5818_ = new_n4835_ & new_n264_;
  assign new_n5819_ = ~new_n5818_;
  assign new_n5820_ = new_n4821_ & shift6;
  assign new_n5821_ = ~new_n5820_;
  assign new_n5822_ = new_n5821_ & new_n5819_;
  assign ores102 = ~new_n5822_;
  assign new_n5824_ = new_n4865_ & new_n264_;
  assign new_n5825_ = ~new_n5824_;
  assign new_n5826_ = new_n4851_ & shift6;
  assign new_n5827_ = ~new_n5826_;
  assign new_n5828_ = new_n5827_ & new_n5825_;
  assign ores103 = ~new_n5828_;
  assign new_n5830_ = new_n4895_ & new_n264_;
  assign new_n5831_ = ~new_n5830_;
  assign new_n5832_ = new_n4881_ & shift6;
  assign new_n5833_ = ~new_n5832_;
  assign new_n5834_ = new_n5833_ & new_n5831_;
  assign ores104 = ~new_n5834_;
  assign new_n5836_ = new_n4925_ & new_n264_;
  assign new_n5837_ = ~new_n5836_;
  assign new_n5838_ = new_n4911_ & shift6;
  assign new_n5839_ = ~new_n5838_;
  assign new_n5840_ = new_n5839_ & new_n5837_;
  assign ores105 = ~new_n5840_;
  assign new_n5842_ = new_n4955_ & new_n264_;
  assign new_n5843_ = ~new_n5842_;
  assign new_n5844_ = new_n4941_ & shift6;
  assign new_n5845_ = ~new_n5844_;
  assign new_n5846_ = new_n5845_ & new_n5843_;
  assign ores106 = ~new_n5846_;
  assign new_n5848_ = new_n4985_ & new_n264_;
  assign new_n5849_ = ~new_n5848_;
  assign new_n5850_ = new_n4971_ & shift6;
  assign new_n5851_ = ~new_n5850_;
  assign new_n5852_ = new_n5851_ & new_n5849_;
  assign ores107 = ~new_n5852_;
  assign new_n5854_ = new_n5015_ & new_n264_;
  assign new_n5855_ = ~new_n5854_;
  assign new_n5856_ = new_n5001_ & shift6;
  assign new_n5857_ = ~new_n5856_;
  assign new_n5858_ = new_n5857_ & new_n5855_;
  assign ores108 = ~new_n5858_;
  assign new_n5860_ = new_n5045_ & new_n264_;
  assign new_n5861_ = ~new_n5860_;
  assign new_n5862_ = new_n5031_ & shift6;
  assign new_n5863_ = ~new_n5862_;
  assign new_n5864_ = new_n5863_ & new_n5861_;
  assign ores109 = ~new_n5864_;
  assign new_n5866_ = new_n5075_ & new_n264_;
  assign new_n5867_ = ~new_n5866_;
  assign new_n5868_ = new_n5061_ & shift6;
  assign new_n5869_ = ~new_n5868_;
  assign new_n5870_ = new_n5869_ & new_n5867_;
  assign ores110 = ~new_n5870_;
  assign new_n5872_ = new_n5105_ & new_n264_;
  assign new_n5873_ = ~new_n5872_;
  assign new_n5874_ = new_n5091_ & shift6;
  assign new_n5875_ = ~new_n5874_;
  assign new_n5876_ = new_n5875_ & new_n5873_;
  assign ores111 = ~new_n5876_;
  assign new_n5878_ = new_n5135_ & new_n264_;
  assign new_n5879_ = ~new_n5878_;
  assign new_n5880_ = new_n5121_ & shift6;
  assign new_n5881_ = ~new_n5880_;
  assign new_n5882_ = new_n5881_ & new_n5879_;
  assign ores112 = ~new_n5882_;
  assign new_n5884_ = new_n5165_ & new_n264_;
  assign new_n5885_ = ~new_n5884_;
  assign new_n5886_ = new_n5151_ & shift6;
  assign new_n5887_ = ~new_n5886_;
  assign new_n5888_ = new_n5887_ & new_n5885_;
  assign ores113 = ~new_n5888_;
  assign new_n5890_ = new_n5195_ & new_n264_;
  assign new_n5891_ = ~new_n5890_;
  assign new_n5892_ = new_n5181_ & shift6;
  assign new_n5893_ = ~new_n5892_;
  assign new_n5894_ = new_n5893_ & new_n5891_;
  assign ores114 = ~new_n5894_;
  assign new_n5896_ = new_n5225_ & new_n264_;
  assign new_n5897_ = ~new_n5896_;
  assign new_n5898_ = new_n5211_ & shift6;
  assign new_n5899_ = ~new_n5898_;
  assign new_n5900_ = new_n5899_ & new_n5897_;
  assign ores115 = ~new_n5900_;
  assign new_n5902_ = new_n5255_ & new_n264_;
  assign new_n5903_ = ~new_n5902_;
  assign new_n5904_ = new_n5241_ & shift6;
  assign new_n5905_ = ~new_n5904_;
  assign new_n5906_ = new_n5905_ & new_n5903_;
  assign ores116 = ~new_n5906_;
  assign new_n5908_ = new_n5285_ & new_n264_;
  assign new_n5909_ = ~new_n5908_;
  assign new_n5910_ = new_n5271_ & shift6;
  assign new_n5911_ = ~new_n5910_;
  assign new_n5912_ = new_n5911_ & new_n5909_;
  assign ores117 = ~new_n5912_;
  assign new_n5914_ = new_n5315_ & new_n264_;
  assign new_n5915_ = ~new_n5914_;
  assign new_n5916_ = new_n5301_ & shift6;
  assign new_n5917_ = ~new_n5916_;
  assign new_n5918_ = new_n5917_ & new_n5915_;
  assign ores118 = ~new_n5918_;
  assign new_n5920_ = new_n5345_ & new_n264_;
  assign new_n5921_ = ~new_n5920_;
  assign new_n5922_ = new_n5331_ & shift6;
  assign new_n5923_ = ~new_n5922_;
  assign new_n5924_ = new_n5923_ & new_n5921_;
  assign ores119 = ~new_n5924_;
  assign new_n5926_ = new_n5375_ & new_n264_;
  assign new_n5927_ = ~new_n5926_;
  assign new_n5928_ = new_n5361_ & shift6;
  assign new_n5929_ = ~new_n5928_;
  assign new_n5930_ = new_n5929_ & new_n5927_;
  assign ores120 = ~new_n5930_;
  assign new_n5932_ = new_n5405_ & new_n264_;
  assign new_n5933_ = ~new_n5932_;
  assign new_n5934_ = new_n5391_ & shift6;
  assign new_n5935_ = ~new_n5934_;
  assign new_n5936_ = new_n5935_ & new_n5933_;
  assign ores121 = ~new_n5936_;
  assign new_n5938_ = new_n5435_ & new_n264_;
  assign new_n5939_ = ~new_n5938_;
  assign new_n5940_ = new_n5421_ & shift6;
  assign new_n5941_ = ~new_n5940_;
  assign new_n5942_ = new_n5941_ & new_n5939_;
  assign ores122 = ~new_n5942_;
  assign new_n5944_ = new_n5465_ & new_n264_;
  assign new_n5945_ = ~new_n5944_;
  assign new_n5946_ = new_n5451_ & shift6;
  assign new_n5947_ = ~new_n5946_;
  assign new_n5948_ = new_n5947_ & new_n5945_;
  assign ores123 = ~new_n5948_;
  assign new_n5950_ = new_n5495_ & new_n264_;
  assign new_n5951_ = ~new_n5950_;
  assign new_n5952_ = new_n5481_ & shift6;
  assign new_n5953_ = ~new_n5952_;
  assign new_n5954_ = new_n5953_ & new_n5951_;
  assign ores124 = ~new_n5954_;
  assign new_n5956_ = new_n5525_ & new_n264_;
  assign new_n5957_ = ~new_n5956_;
  assign new_n5958_ = new_n5511_ & shift6;
  assign new_n5959_ = ~new_n5958_;
  assign new_n5960_ = new_n5959_ & new_n5957_;
  assign ores125 = ~new_n5960_;
  assign new_n5962_ = new_n5555_ & new_n264_;
  assign new_n5963_ = ~new_n5962_;
  assign new_n5964_ = new_n5541_ & shift6;
  assign new_n5965_ = ~new_n5964_;
  assign new_n5966_ = new_n5965_ & new_n5963_;
  assign ores126 = ~new_n5966_;
  assign new_n5968_ = new_n5585_ & new_n264_;
  assign new_n5969_ = ~new_n5968_;
  assign new_n5970_ = new_n5571_ & shift6;
  assign new_n5971_ = ~new_n5970_;
  assign new_n5972_ = new_n5971_ & new_n5969_;
  assign ores127 = ~new_n5972_;
endmodule


