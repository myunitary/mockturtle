// Benchmark "/tmp/tmp" written by ABC on Wed Nov 12 17:56:38 2025

module FP-eq_opt ( 
    n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
    n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63  );
  input  n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
    n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9, po10, po11, po12,
    po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24,
    po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36,
    po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48,
    po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60,
    po61, po62, po63;
  wire new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582;
  assign new_n129 = n61 & n62;
  assign new_n130 = n63 & new_n129;
  assign new_n131 = n53 & n54;
  assign new_n132 = n55 & n56;
  assign new_n133 = new_n131 & new_n132;
  assign new_n134 = n59 & n60;
  assign new_n135 = n57 & n58;
  assign new_n136 = new_n134 & new_n135;
  assign new_n137 = new_n133 & new_n136;
  assign new_n138 = new_n130 & new_n137;
  assign new_n139 = ~n51 & ~n52;
  assign new_n140 = ~n49 & ~n50;
  assign new_n141 = new_n139 & new_n140;
  assign new_n142 = ~n47 & ~n48;
  assign new_n143 = ~n45 & ~n46;
  assign new_n144 = new_n142 & new_n143;
  assign new_n145 = ~n43 & ~n44;
  assign new_n146 = ~n41 & ~n42;
  assign new_n147 = new_n145 & new_n146;
  assign new_n148 = new_n144 & new_n147;
  assign new_n149 = ~n39 & ~n40;
  assign new_n150 = ~n37 & ~n38;
  assign new_n151 = new_n149 & new_n150;
  assign new_n152 = ~n35 & ~n36;
  assign new_n153 = ~n33 & ~n34;
  assign new_n154 = new_n152 & new_n153;
  assign new_n155 = new_n151 & new_n154;
  assign new_n156 = new_n148 & new_n155;
  assign new_n157 = new_n141 & new_n156;
  assign new_n158 = ~n31 & ~n32;
  assign new_n159 = ~n29 & ~n30;
  assign new_n160 = new_n158 & new_n159;
  assign new_n161 = ~n27 & ~n28;
  assign new_n162 = ~n25 & ~n26;
  assign new_n163 = new_n161 & new_n162;
  assign new_n164 = new_n160 & new_n163;
  assign new_n165 = ~n23 & ~n24;
  assign new_n166 = ~n21 & ~n22;
  assign new_n167 = new_n165 & new_n166;
  assign new_n168 = ~n19 & ~n20;
  assign new_n169 = ~n17 & ~n18;
  assign new_n170 = new_n168 & new_n169;
  assign new_n171 = new_n167 & new_n170;
  assign new_n172 = new_n164 & new_n171;
  assign new_n173 = ~n15 & ~n16;
  assign new_n174 = ~n13 & ~n14;
  assign new_n175 = new_n173 & new_n174;
  assign new_n176 = ~n11 & ~n12;
  assign new_n177 = ~n9 & ~n10;
  assign new_n178 = new_n176 & new_n177;
  assign new_n179 = new_n175 & new_n178;
  assign new_n180 = ~n7 & ~n8;
  assign new_n181 = ~n5 & ~n6;
  assign new_n182 = new_n180 & new_n181;
  assign new_n183 = ~n3 & ~n4;
  assign new_n184 = ~n1 & ~n2;
  assign new_n185 = new_n183 & new_n184;
  assign new_n186 = new_n182 & new_n185;
  assign new_n187 = new_n179 & new_n186;
  assign new_n188 = new_n172 & new_n187;
  assign new_n189 = new_n157 & new_n188;
  assign new_n190 = ~new_n189 & new_n138;
  assign new_n191 = n125 & n126;
  assign new_n192 = n127 & new_n191;
  assign new_n193 = n123 & n124;
  assign new_n194 = n121 & n122;
  assign new_n195 = new_n193 & new_n194;
  assign new_n196 = n117 & n118;
  assign new_n197 = n119 & n120;
  assign new_n198 = new_n196 & new_n197;
  assign new_n199 = new_n195 & new_n198;
  assign new_n200 = new_n192 & new_n199;
  assign new_n201 = ~n115 & ~n116;
  assign new_n202 = ~n113 & ~n114;
  assign new_n203 = new_n201 & new_n202;
  assign new_n204 = ~n111 & ~n112;
  assign new_n205 = ~n109 & ~n110;
  assign new_n206 = new_n204 & new_n205;
  assign new_n207 = ~n107 & ~n108;
  assign new_n208 = ~n105 & ~n106;
  assign new_n209 = new_n207 & new_n208;
  assign new_n210 = new_n206 & new_n209;
  assign new_n211 = ~n103 & ~n104;
  assign new_n212 = ~n101 & ~n102;
  assign new_n213 = new_n211 & new_n212;
  assign new_n214 = ~n99 & ~n100;
  assign new_n215 = ~n97 & ~n98;
  assign new_n216 = new_n214 & new_n215;
  assign new_n217 = new_n213 & new_n216;
  assign new_n218 = new_n210 & new_n217;
  assign new_n219 = new_n203 & new_n218;
  assign new_n220 = ~n95 & ~n96;
  assign new_n221 = ~n93 & ~n94;
  assign new_n222 = new_n220 & new_n221;
  assign new_n223 = ~n91 & ~n92;
  assign new_n224 = ~n89 & ~n90;
  assign new_n225 = new_n223 & new_n224;
  assign new_n226 = new_n222 & new_n225;
  assign new_n227 = ~n87 & ~n88;
  assign new_n228 = ~n85 & ~n86;
  assign new_n229 = new_n227 & new_n228;
  assign new_n230 = ~n83 & ~n84;
  assign new_n231 = ~n81 & ~n82;
  assign new_n232 = new_n230 & new_n231;
  assign new_n233 = new_n229 & new_n232;
  assign new_n234 = new_n226 & new_n233;
  assign new_n235 = ~n79 & ~n80;
  assign new_n236 = ~n77 & ~n78;
  assign new_n237 = new_n235 & new_n236;
  assign new_n238 = ~n75 & ~n76;
  assign new_n239 = ~n73 & ~n74;
  assign new_n240 = new_n238 & new_n239;
  assign new_n241 = new_n237 & new_n240;
  assign new_n242 = ~n71 & ~n72;
  assign new_n243 = ~n69 & ~n70;
  assign new_n244 = new_n242 & new_n243;
  assign new_n245 = ~n67 & ~n68;
  assign new_n246 = ~n65 & ~n66;
  assign new_n247 = new_n245 & new_n246;
  assign new_n248 = new_n244 & new_n247;
  assign new_n249 = new_n241 & new_n248;
  assign new_n250 = new_n234 & new_n249;
  assign new_n251 = new_n219 & new_n250;
  assign new_n252 = ~new_n251 & new_n200;
  assign new_n253 = ~new_n190 & ~new_n252;
  assign new_n254 = n127 ^ n124;
  assign new_n255 = ~n125 & new_n254;
  assign new_n256 = new_n255 ^ n125;
  assign new_n257 = new_n255 ^ n126;
  assign new_n258 = ~n127 & ~new_n257;
  assign new_n259 = new_n258 ^ n127;
  assign new_n260 = new_n259 ^ n124;
  assign new_n261 = ~new_n256 & new_n260;
  assign new_n262 = ~n62 & ~n63;
  assign new_n263 = ~n60 & ~n61;
  assign new_n264 = new_n262 & new_n263;
  assign new_n265 = new_n261 & new_n264;
  assign new_n266 = n123 ^ n120;
  assign new_n267 = ~n121 & new_n266;
  assign new_n268 = new_n267 ^ n121;
  assign new_n269 = new_n267 ^ n122;
  assign new_n270 = ~n123 & ~new_n269;
  assign new_n271 = new_n270 ^ n123;
  assign new_n272 = new_n271 ^ n120;
  assign new_n273 = ~new_n268 & new_n272;
  assign new_n274 = ~n58 & ~n59;
  assign new_n275 = ~n56 & ~n57;
  assign new_n276 = new_n274 & new_n275;
  assign new_n277 = new_n273 & new_n276;
  assign new_n278 = new_n265 & new_n277;
  assign new_n279 = n119 ^ n116;
  assign new_n280 = ~n117 & new_n279;
  assign new_n281 = new_n280 ^ n117;
  assign new_n282 = new_n280 ^ n118;
  assign new_n283 = ~n119 & ~new_n282;
  assign new_n284 = new_n283 ^ n119;
  assign new_n285 = new_n284 ^ n116;
  assign new_n286 = ~new_n281 & new_n285;
  assign new_n287 = ~n54 & ~n55;
  assign new_n288 = ~n52 & ~n53;
  assign new_n289 = new_n287 & new_n288;
  assign new_n290 = new_n286 & new_n289;
  assign new_n291 = n115 ^ n112;
  assign new_n292 = ~n113 & new_n291;
  assign new_n293 = new_n292 ^ n113;
  assign new_n294 = new_n292 ^ n114;
  assign new_n295 = ~n115 & ~new_n294;
  assign new_n296 = new_n295 ^ n115;
  assign new_n297 = new_n296 ^ n112;
  assign new_n298 = ~new_n293 & new_n297;
  assign new_n299 = ~n50 & ~n51;
  assign new_n300 = ~n48 & ~n49;
  assign new_n301 = new_n299 & new_n300;
  assign new_n302 = new_n298 & new_n301;
  assign new_n303 = new_n290 & new_n302;
  assign new_n304 = new_n278 & new_n303;
  assign new_n305 = n111 ^ n108;
  assign new_n306 = ~n109 & new_n305;
  assign new_n307 = new_n306 ^ n109;
  assign new_n308 = new_n306 ^ n110;
  assign new_n309 = ~n111 & ~new_n308;
  assign new_n310 = new_n309 ^ n111;
  assign new_n311 = new_n310 ^ n108;
  assign new_n312 = ~new_n307 & new_n311;
  assign new_n313 = ~n46 & ~n47;
  assign new_n314 = ~n44 & ~n45;
  assign new_n315 = new_n313 & new_n314;
  assign new_n316 = new_n312 & new_n315;
  assign new_n317 = n107 ^ n104;
  assign new_n318 = ~n105 & new_n317;
  assign new_n319 = new_n318 ^ n105;
  assign new_n320 = new_n318 ^ n106;
  assign new_n321 = ~n107 & ~new_n320;
  assign new_n322 = new_n321 ^ n107;
  assign new_n323 = new_n322 ^ n104;
  assign new_n324 = ~new_n319 & new_n323;
  assign new_n325 = ~n42 & ~n43;
  assign new_n326 = ~n40 & ~n41;
  assign new_n327 = new_n325 & new_n326;
  assign new_n328 = new_n324 & new_n327;
  assign new_n329 = new_n316 & new_n328;
  assign new_n330 = n103 ^ n100;
  assign new_n331 = ~n101 & new_n330;
  assign new_n332 = new_n331 ^ n101;
  assign new_n333 = new_n331 ^ n102;
  assign new_n334 = ~n103 & ~new_n333;
  assign new_n335 = new_n334 ^ n103;
  assign new_n336 = new_n335 ^ n100;
  assign new_n337 = ~new_n332 & new_n336;
  assign new_n338 = ~n38 & ~n39;
  assign new_n339 = ~n36 & ~n37;
  assign new_n340 = new_n338 & new_n339;
  assign new_n341 = new_n337 & new_n340;
  assign new_n342 = n99 ^ n96;
  assign new_n343 = ~n97 & new_n342;
  assign new_n344 = new_n343 ^ n97;
  assign new_n345 = new_n343 ^ n98;
  assign new_n346 = ~n99 & ~new_n345;
  assign new_n347 = new_n346 ^ n99;
  assign new_n348 = new_n347 ^ n96;
  assign new_n349 = ~new_n344 & new_n348;
  assign new_n350 = ~n34 & ~n35;
  assign new_n351 = ~n32 & ~n33;
  assign new_n352 = new_n350 & new_n351;
  assign new_n353 = new_n349 & new_n352;
  assign new_n354 = new_n341 & new_n353;
  assign new_n355 = new_n329 & new_n354;
  assign new_n356 = new_n304 & new_n355;
  assign new_n357 = n95 ^ n92;
  assign new_n358 = ~n93 & new_n357;
  assign new_n359 = new_n358 ^ n93;
  assign new_n360 = new_n358 ^ n94;
  assign new_n361 = ~n95 & ~new_n360;
  assign new_n362 = new_n361 ^ n95;
  assign new_n363 = new_n362 ^ n92;
  assign new_n364 = ~new_n359 & new_n363;
  assign new_n365 = ~n30 & ~n31;
  assign new_n366 = ~n28 & ~n29;
  assign new_n367 = new_n365 & new_n366;
  assign new_n368 = new_n364 & new_n367;
  assign new_n369 = n91 ^ n88;
  assign new_n370 = ~n89 & new_n369;
  assign new_n371 = new_n370 ^ n89;
  assign new_n372 = new_n370 ^ n90;
  assign new_n373 = ~n91 & ~new_n372;
  assign new_n374 = new_n373 ^ n91;
  assign new_n375 = new_n374 ^ n88;
  assign new_n376 = ~new_n371 & new_n375;
  assign new_n377 = ~n26 & ~n27;
  assign new_n378 = ~n24 & ~n25;
  assign new_n379 = new_n377 & new_n378;
  assign new_n380 = new_n376 & new_n379;
  assign new_n381 = new_n368 & new_n380;
  assign new_n382 = n87 ^ n84;
  assign new_n383 = ~n85 & new_n382;
  assign new_n384 = new_n383 ^ n85;
  assign new_n385 = new_n383 ^ n86;
  assign new_n386 = ~n87 & ~new_n385;
  assign new_n387 = new_n386 ^ n87;
  assign new_n388 = new_n387 ^ n84;
  assign new_n389 = ~new_n384 & new_n388;
  assign new_n390 = ~n22 & ~n23;
  assign new_n391 = ~n20 & ~n21;
  assign new_n392 = new_n390 & new_n391;
  assign new_n393 = new_n389 & new_n392;
  assign new_n394 = n83 ^ n80;
  assign new_n395 = ~n81 & new_n394;
  assign new_n396 = new_n395 ^ n81;
  assign new_n397 = new_n395 ^ n82;
  assign new_n398 = ~n83 & ~new_n397;
  assign new_n399 = new_n398 ^ n83;
  assign new_n400 = new_n399 ^ n80;
  assign new_n401 = ~new_n396 & new_n400;
  assign new_n402 = ~n18 & ~n19;
  assign new_n403 = ~n16 & ~n17;
  assign new_n404 = new_n402 & new_n403;
  assign new_n405 = new_n401 & new_n404;
  assign new_n406 = new_n393 & new_n405;
  assign new_n407 = new_n381 & new_n406;
  assign new_n408 = n79 ^ n76;
  assign new_n409 = ~n77 & new_n408;
  assign new_n410 = new_n409 ^ n77;
  assign new_n411 = new_n409 ^ n78;
  assign new_n412 = ~n79 & ~new_n411;
  assign new_n413 = new_n412 ^ n79;
  assign new_n414 = new_n413 ^ n76;
  assign new_n415 = ~new_n410 & new_n414;
  assign new_n416 = ~n14 & ~n15;
  assign new_n417 = ~n12 & ~n13;
  assign new_n418 = new_n416 & new_n417;
  assign new_n419 = new_n415 & new_n418;
  assign new_n420 = n75 ^ n72;
  assign new_n421 = ~n73 & new_n420;
  assign new_n422 = new_n421 ^ n73;
  assign new_n423 = new_n421 ^ n74;
  assign new_n424 = ~n75 & ~new_n423;
  assign new_n425 = new_n424 ^ n75;
  assign new_n426 = new_n425 ^ n72;
  assign new_n427 = ~new_n422 & new_n426;
  assign new_n428 = ~n10 & ~n11;
  assign new_n429 = ~n8 & ~n9;
  assign new_n430 = new_n428 & new_n429;
  assign new_n431 = new_n427 & new_n430;
  assign new_n432 = new_n419 & new_n431;
  assign new_n433 = ~n66 & ~n67;
  assign new_n434 = ~n65 & new_n433;
  assign new_n435 = ~n2 & ~n3;
  assign new_n436 = ~n1 & new_n435;
  assign new_n437 = new_n434 & new_n436;
  assign new_n438 = n71 ^ n68;
  assign new_n439 = ~n69 & new_n438;
  assign new_n440 = new_n439 ^ n69;
  assign new_n441 = new_n439 ^ n70;
  assign new_n442 = ~n71 & ~new_n441;
  assign new_n443 = new_n442 ^ n71;
  assign new_n444 = new_n443 ^ n68;
  assign new_n445 = ~new_n440 & new_n444;
  assign new_n446 = ~n6 & ~n7;
  assign new_n447 = ~n4 & ~n5;
  assign new_n448 = new_n446 & new_n447;
  assign new_n449 = new_n445 & new_n448;
  assign new_n450 = new_n437 & new_n449;
  assign new_n451 = new_n432 & new_n450;
  assign new_n452 = new_n407 & new_n451;
  assign new_n453 = new_n356 & new_n452;
  assign new_n454 = n128 ^ n64;
  assign new_n455 = n127 ^ n63;
  assign new_n456 = ~new_n454 & ~new_n455;
  assign new_n457 = n126 ^ n62;
  assign new_n458 = n125 ^ n61;
  assign new_n459 = ~new_n457 & ~new_n458;
  assign new_n460 = new_n456 & new_n459;
  assign new_n461 = n124 ^ n60;
  assign new_n462 = n123 ^ n59;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = n122 ^ n58;
  assign new_n465 = n121 ^ n57;
  assign new_n466 = ~new_n464 & ~new_n465;
  assign new_n467 = new_n463 & new_n466;
  assign new_n468 = new_n460 & new_n467;
  assign new_n469 = n120 ^ n56;
  assign new_n470 = n119 ^ n55;
  assign new_n471 = ~new_n469 & ~new_n470;
  assign new_n472 = n118 ^ n54;
  assign new_n473 = n117 ^ n53;
  assign new_n474 = ~new_n472 & ~new_n473;
  assign new_n475 = new_n471 & new_n474;
  assign new_n476 = n116 ^ n52;
  assign new_n477 = n115 ^ n51;
  assign new_n478 = ~new_n476 & ~new_n477;
  assign new_n479 = n114 ^ n50;
  assign new_n480 = n113 ^ n49;
  assign new_n481 = ~new_n479 & ~new_n480;
  assign new_n482 = new_n478 & new_n481;
  assign new_n483 = new_n475 & new_n482;
  assign new_n484 = new_n468 & new_n483;
  assign new_n485 = n112 ^ n48;
  assign new_n486 = n111 ^ n47;
  assign new_n487 = ~new_n485 & ~new_n486;
  assign new_n488 = n110 ^ n46;
  assign new_n489 = n109 ^ n45;
  assign new_n490 = ~new_n488 & ~new_n489;
  assign new_n491 = new_n487 & new_n490;
  assign new_n492 = n108 ^ n44;
  assign new_n493 = n107 ^ n43;
  assign new_n494 = ~new_n492 & ~new_n493;
  assign new_n495 = n106 ^ n42;
  assign new_n496 = n105 ^ n41;
  assign new_n497 = ~new_n495 & ~new_n496;
  assign new_n498 = new_n494 & new_n497;
  assign new_n499 = new_n491 & new_n498;
  assign new_n500 = n104 ^ n40;
  assign new_n501 = n103 ^ n39;
  assign new_n502 = ~new_n500 & ~new_n501;
  assign new_n503 = n102 ^ n38;
  assign new_n504 = n101 ^ n37;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = new_n502 & new_n505;
  assign new_n507 = n100 ^ n36;
  assign new_n508 = n99 ^ n35;
  assign new_n509 = ~new_n507 & ~new_n508;
  assign new_n510 = n98 ^ n34;
  assign new_n511 = n97 ^ n33;
  assign new_n512 = ~new_n510 & ~new_n511;
  assign new_n513 = new_n509 & new_n512;
  assign new_n514 = new_n506 & new_n513;
  assign new_n515 = new_n499 & new_n514;
  assign new_n516 = new_n484 & new_n515;
  assign new_n517 = n96 ^ n32;
  assign new_n518 = n95 ^ n31;
  assign new_n519 = ~new_n517 & ~new_n518;
  assign new_n520 = n94 ^ n30;
  assign new_n521 = n93 ^ n29;
  assign new_n522 = ~new_n520 & ~new_n521;
  assign new_n523 = new_n519 & new_n522;
  assign new_n524 = n92 ^ n28;
  assign new_n525 = n91 ^ n27;
  assign new_n526 = ~new_n524 & ~new_n525;
  assign new_n527 = n90 ^ n26;
  assign new_n528 = n89 ^ n25;
  assign new_n529 = ~new_n527 & ~new_n528;
  assign new_n530 = new_n526 & new_n529;
  assign new_n531 = new_n523 & new_n530;
  assign new_n532 = n88 ^ n24;
  assign new_n533 = n87 ^ n23;
  assign new_n534 = ~new_n532 & ~new_n533;
  assign new_n535 = n86 ^ n22;
  assign new_n536 = n85 ^ n21;
  assign new_n537 = ~new_n535 & ~new_n536;
  assign new_n538 = new_n534 & new_n537;
  assign new_n539 = n84 ^ n20;
  assign new_n540 = n83 ^ n19;
  assign new_n541 = ~new_n539 & ~new_n540;
  assign new_n542 = n82 ^ n18;
  assign new_n543 = n81 ^ n17;
  assign new_n544 = ~new_n542 & ~new_n543;
  assign new_n545 = new_n541 & new_n544;
  assign new_n546 = new_n538 & new_n545;
  assign new_n547 = new_n531 & new_n546;
  assign new_n548 = n80 ^ n16;
  assign new_n549 = n79 ^ n15;
  assign new_n550 = ~new_n548 & ~new_n549;
  assign new_n551 = n78 ^ n14;
  assign new_n552 = n77 ^ n13;
  assign new_n553 = ~new_n551 & ~new_n552;
  assign new_n554 = new_n550 & new_n553;
  assign new_n555 = n76 ^ n12;
  assign new_n556 = n75 ^ n11;
  assign new_n557 = ~new_n555 & ~new_n556;
  assign new_n558 = n74 ^ n10;
  assign new_n559 = n73 ^ n9;
  assign new_n560 = ~new_n558 & ~new_n559;
  assign new_n561 = new_n557 & new_n560;
  assign new_n562 = new_n554 & new_n561;
  assign new_n563 = n72 ^ n8;
  assign new_n564 = n71 ^ n7;
  assign new_n565 = ~new_n563 & ~new_n564;
  assign new_n566 = n70 ^ n6;
  assign new_n567 = n69 ^ n5;
  assign new_n568 = ~new_n566 & ~new_n567;
  assign new_n569 = new_n565 & new_n568;
  assign new_n570 = n68 ^ n4;
  assign new_n571 = n67 ^ n3;
  assign new_n572 = ~new_n570 & ~new_n571;
  assign new_n573 = n66 ^ n2;
  assign new_n574 = n65 ^ n1;
  assign new_n575 = ~new_n573 & ~new_n574;
  assign new_n576 = new_n572 & new_n575;
  assign new_n577 = new_n569 & new_n576;
  assign new_n578 = new_n562 & new_n577;
  assign new_n579 = new_n547 & new_n578;
  assign new_n580 = new_n516 & new_n579;
  assign new_n581 = ~new_n453 & ~new_n580;
  assign new_n582 = ~new_n581 & new_n253;
  assign po0 = new_n582;
  assign po1 = 1'b0;
  assign po2 = 1'b0;
  assign po3 = 1'b0;
  assign po4 = 1'b0;
  assign po5 = 1'b0;
  assign po6 = 1'b0;
  assign po7 = 1'b0;
  assign po8 = 1'b0;
  assign po9 = 1'b0;
  assign po10 = 1'b0;
  assign po11 = 1'b0;
  assign po12 = 1'b0;
  assign po13 = 1'b0;
  assign po14 = 1'b0;
  assign po15 = 1'b0;
  assign po16 = 1'b0;
  assign po17 = 1'b0;
  assign po18 = 1'b0;
  assign po19 = 1'b0;
  assign po20 = 1'b0;
  assign po21 = 1'b0;
  assign po22 = 1'b0;
  assign po23 = 1'b0;
  assign po24 = 1'b0;
  assign po25 = 1'b0;
  assign po26 = 1'b0;
  assign po27 = 1'b0;
  assign po28 = 1'b0;
  assign po29 = 1'b0;
  assign po30 = 1'b0;
  assign po31 = 1'b0;
  assign po32 = 1'b0;
  assign po33 = 1'b0;
  assign po34 = 1'b0;
  assign po35 = 1'b0;
  assign po36 = 1'b0;
  assign po37 = 1'b0;
  assign po38 = 1'b0;
  assign po39 = 1'b0;
  assign po40 = 1'b0;
  assign po41 = 1'b0;
  assign po42 = 1'b0;
  assign po43 = 1'b0;
  assign po44 = 1'b0;
  assign po45 = 1'b0;
  assign po46 = 1'b0;
  assign po47 = 1'b0;
  assign po48 = 1'b0;
  assign po49 = 1'b0;
  assign po50 = 1'b0;
  assign po51 = 1'b0;
  assign po52 = 1'b0;
  assign po53 = 1'b0;
  assign po54 = 1'b0;
  assign po55 = 1'b0;
  assign po56 = 1'b0;
  assign po57 = 1'b0;
  assign po58 = 1'b0;
  assign po59 = 1'b0;
  assign po60 = 1'b0;
  assign po61 = 1'b0;
  assign po62 = 1'b0;
  assign po63 = 1'b0;
endmodule


