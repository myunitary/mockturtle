module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 ;
  wire n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 ;
  assign n289 = ~x94 & ~x286 ;
  assign n290 = x94 & x286 ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = ~x93 & ~x285 ;
  assign n293 = x93 & x285 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = n291 & n294 ;
  assign n296 = ~n291 & ~n294 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = ~x95 & ~x287 ;
  assign n299 = x95 & x287 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = ~n297 & ~n300 ;
  assign n302 = n297 & n300 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~x89 & ~x281 ;
  assign n305 = x89 & x281 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = ~n303 & ~n306 ;
  assign n308 = n303 & n306 ;
  assign n309 = ~n307 & ~n308 ;
  assign n310 = ~x91 & ~x283 ;
  assign n311 = x91 & x283 ;
  assign n312 = ~n310 & ~n311 ;
  assign n313 = ~x90 & ~x282 ;
  assign n314 = x90 & x282 ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = ~n312 & ~n315 ;
  assign n317 = n312 & n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~x92 & ~x284 ;
  assign n320 = x92 & x284 ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = ~n318 & ~n321 ;
  assign n323 = n318 & n321 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n309 & ~n324 ;
  assign n326 = ~n307 & ~n325 ;
  assign n327 = ~n295 & ~n302 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = n326 & ~n327 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n317 & ~n323 ;
  assign n332 = n330 & n331 ;
  assign n333 = ~n328 & ~n332 ;
  assign n334 = ~n330 & ~n331 ;
  assign n335 = ~n332 & ~n334 ;
  assign n336 = ~n309 & n324 ;
  assign n337 = ~n325 & ~n336 ;
  assign n338 = ~x81 & ~x273 ;
  assign n339 = x81 & x273 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n337 & ~n340 ;
  assign n342 = ~x87 & ~x279 ;
  assign n343 = x87 & x279 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = ~x86 & ~x278 ;
  assign n346 = x86 & x278 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n344 & ~n347 ;
  assign n349 = n344 & n347 ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = ~x88 & ~x280 ;
  assign n352 = x88 & x280 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = ~n350 & ~n353 ;
  assign n355 = n350 & n353 ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = ~x82 & ~x274 ;
  assign n358 = x82 & x274 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = ~n356 & ~n359 ;
  assign n361 = n356 & n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~x84 & ~x276 ;
  assign n364 = x84 & x276 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = ~x83 & ~x275 ;
  assign n367 = x83 & x275 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = ~n365 & ~n368 ;
  assign n370 = n365 & n368 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = ~x85 & ~x277 ;
  assign n373 = x85 & x277 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = ~n371 & ~n374 ;
  assign n376 = n371 & n374 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = n362 & ~n377 ;
  assign n379 = ~n362 & n377 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n337 & n340 ;
  assign n382 = ~n341 & ~n381 ;
  assign n383 = n380 & n382 ;
  assign n384 = ~n341 & ~n383 ;
  assign n385 = n335 & ~n384 ;
  assign n386 = ~n360 & ~n378 ;
  assign n387 = ~n349 & ~n355 ;
  assign n388 = ~n386 & n387 ;
  assign n389 = n386 & ~n387 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = ~n370 & ~n376 ;
  assign n392 = n390 & n391 ;
  assign n393 = ~n390 & ~n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n335 & n384 ;
  assign n396 = ~n385 & ~n395 ;
  assign n397 = n394 & n396 ;
  assign n398 = ~n385 & ~n397 ;
  assign n399 = ~n333 & ~n398 ;
  assign n400 = n333 & n398 ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = ~n388 & ~n392 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = ~n399 & ~n403 ;
  assign n405 = ~n401 & n402 ;
  assign n406 = ~n403 & ~n405 ;
  assign n407 = ~n394 & ~n396 ;
  assign n408 = ~n397 & ~n407 ;
  assign n409 = ~n380 & ~n382 ;
  assign n410 = ~n383 & ~n409 ;
  assign n411 = ~x65 & ~x257 ;
  assign n412 = x65 & x257 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = n410 & ~n413 ;
  assign n415 = ~x72 & ~x264 ;
  assign n416 = x72 & x264 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = ~x71 & ~x263 ;
  assign n419 = x71 & x263 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n417 & ~n420 ;
  assign n422 = n417 & n420 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~x73 & ~x265 ;
  assign n425 = x73 & x265 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~n423 & ~n426 ;
  assign n428 = n423 & n426 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = ~x67 & ~x259 ;
  assign n431 = x67 & x259 ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = ~n429 & ~n432 ;
  assign n434 = n429 & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = ~x69 & ~x261 ;
  assign n437 = x69 & x261 ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = ~x68 & ~x260 ;
  assign n440 = x68 & x260 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~n438 & ~n441 ;
  assign n443 = n438 & n441 ;
  assign n444 = ~n442 & ~n443 ;
  assign n445 = ~x70 & ~x262 ;
  assign n446 = x70 & x262 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n444 & ~n447 ;
  assign n449 = n444 & n447 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = n435 & ~n450 ;
  assign n452 = ~n435 & n450 ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = ~x79 & ~x271 ;
  assign n455 = x79 & x271 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = ~x78 & ~x270 ;
  assign n458 = x78 & x270 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = ~n456 & ~n459 ;
  assign n461 = n456 & n459 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~x80 & ~x272 ;
  assign n464 = x80 & x272 ;
  assign n465 = ~n463 & ~n464 ;
  assign n466 = ~n462 & ~n465 ;
  assign n467 = n462 & n465 ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = ~x74 & ~x266 ;
  assign n470 = x74 & x266 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~n468 & ~n471 ;
  assign n473 = n468 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~x76 & ~x268 ;
  assign n476 = x76 & x268 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~x75 & ~x267 ;
  assign n479 = x75 & x267 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = ~n477 & ~n480 ;
  assign n482 = n477 & n480 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = ~x77 & ~x269 ;
  assign n485 = x77 & x269 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~n483 & ~n486 ;
  assign n488 = n483 & n486 ;
  assign n489 = ~n487 & ~n488 ;
  assign n490 = n474 & ~n489 ;
  assign n491 = ~n474 & n489 ;
  assign n492 = ~n490 & ~n491 ;
  assign n493 = ~x66 & ~x258 ;
  assign n494 = x66 & x258 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n492 & ~n495 ;
  assign n497 = ~n492 & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = n453 & n498 ;
  assign n500 = ~n453 & ~n498 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = ~n410 & n413 ;
  assign n503 = ~n414 & ~n502 ;
  assign n504 = n501 & n503 ;
  assign n505 = ~n414 & ~n504 ;
  assign n506 = n408 & ~n505 ;
  assign n507 = ~n433 & ~n451 ;
  assign n508 = ~n422 & ~n428 ;
  assign n509 = ~n507 & n508 ;
  assign n510 = n507 & ~n508 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = ~n443 & ~n449 ;
  assign n513 = n511 & n512 ;
  assign n514 = ~n511 & ~n512 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = ~n472 & ~n490 ;
  assign n517 = ~n461 & ~n467 ;
  assign n518 = ~n516 & n517 ;
  assign n519 = n516 & ~n517 ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = ~n482 & ~n488 ;
  assign n522 = n520 & n521 ;
  assign n523 = ~n520 & ~n521 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n496 & ~n499 ;
  assign n526 = n524 & ~n525 ;
  assign n527 = ~n524 & n525 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = n515 & n528 ;
  assign n530 = ~n515 & ~n528 ;
  assign n531 = ~n529 & ~n530 ;
  assign n532 = ~n408 & n505 ;
  assign n533 = ~n506 & ~n532 ;
  assign n534 = n531 & n533 ;
  assign n535 = ~n506 & ~n534 ;
  assign n536 = n406 & ~n535 ;
  assign n537 = ~n518 & ~n522 ;
  assign n538 = ~n526 & ~n529 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = n537 & n538 ;
  assign n541 = ~n539 & ~n540 ;
  assign n542 = ~n509 & ~n513 ;
  assign n543 = n541 & ~n542 ;
  assign n544 = ~n541 & n542 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~n406 & n535 ;
  assign n547 = ~n536 & ~n546 ;
  assign n548 = n545 & n547 ;
  assign n549 = ~n536 & ~n548 ;
  assign n550 = ~n404 & ~n549 ;
  assign n551 = n404 & n549 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = ~n539 & ~n543 ;
  assign n554 = n552 & ~n553 ;
  assign n555 = ~n550 & ~n554 ;
  assign n556 = ~n552 & n553 ;
  assign n557 = ~n554 & ~n556 ;
  assign n558 = ~n545 & ~n547 ;
  assign n559 = ~n548 & ~n558 ;
  assign n560 = ~n531 & ~n533 ;
  assign n561 = ~n534 & ~n560 ;
  assign n562 = ~n501 & ~n503 ;
  assign n563 = ~n504 & ~n562 ;
  assign n564 = ~x64 & ~x256 ;
  assign n565 = x64 & x256 ;
  assign n566 = ~n564 & ~n565 ;
  assign n567 = ~n563 & n566 ;
  assign n568 = ~n561 & n567 ;
  assign n569 = ~n559 & n568 ;
  assign n570 = ~n557 & n569 ;
  assign n571 = n555 & n570 ;
  assign n572 = ~x254 & ~x286 ;
  assign n573 = x254 & x286 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = ~x253 & ~x285 ;
  assign n576 = x253 & x285 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = n574 & n577 ;
  assign n579 = ~n574 & ~n577 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = ~x255 & ~x287 ;
  assign n582 = x255 & x287 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n580 & n583 ;
  assign n585 = ~n578 & ~n584 ;
  assign n586 = ~n580 & ~n583 ;
  assign n587 = ~n584 & ~n586 ;
  assign n588 = ~x249 & ~x281 ;
  assign n589 = x249 & x281 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = n587 & n590 ;
  assign n592 = ~n587 & ~n590 ;
  assign n593 = ~x251 & ~x283 ;
  assign n594 = x251 & x283 ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = ~x250 & ~x282 ;
  assign n597 = x250 & x282 ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = ~n595 & ~n598 ;
  assign n600 = n595 & n598 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~x252 & ~x284 ;
  assign n603 = x252 & x284 ;
  assign n604 = ~n602 & ~n603 ;
  assign n605 = ~n601 & ~n604 ;
  assign n606 = n601 & n604 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = ~n592 & n607 ;
  assign n609 = ~n591 & ~n608 ;
  assign n610 = n585 & n609 ;
  assign n611 = ~n585 & ~n609 ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = ~n600 & ~n606 ;
  assign n614 = n612 & n613 ;
  assign n615 = ~n610 & ~n614 ;
  assign n616 = ~n612 & ~n613 ;
  assign n617 = ~n614 & ~n616 ;
  assign n618 = ~n591 & ~n592 ;
  assign n619 = ~n607 & n618 ;
  assign n620 = n607 & ~n618 ;
  assign n621 = ~n619 & ~n620 ;
  assign n622 = ~x241 & ~x273 ;
  assign n623 = x241 & x273 ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = ~n621 & n624 ;
  assign n626 = n621 & ~n624 ;
  assign n627 = ~x247 & ~x279 ;
  assign n628 = x247 & x279 ;
  assign n629 = ~n627 & ~n628 ;
  assign n630 = ~x246 & ~x278 ;
  assign n631 = x246 & x278 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = ~n629 & ~n632 ;
  assign n634 = n629 & n632 ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = ~x248 & ~x280 ;
  assign n637 = x248 & x280 ;
  assign n638 = ~n636 & ~n637 ;
  assign n639 = ~n635 & ~n638 ;
  assign n640 = n635 & n638 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = ~x242 & ~x274 ;
  assign n643 = x242 & x274 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = ~n641 & ~n644 ;
  assign n646 = n641 & n644 ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = ~x244 & ~x276 ;
  assign n649 = x244 & x276 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = ~x243 & ~x275 ;
  assign n652 = x243 & x275 ;
  assign n653 = ~n651 & ~n652 ;
  assign n654 = ~n650 & ~n653 ;
  assign n655 = n650 & n653 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~x245 & ~x277 ;
  assign n658 = x245 & x277 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = ~n656 & ~n659 ;
  assign n661 = n656 & n659 ;
  assign n662 = ~n660 & ~n661 ;
  assign n663 = n647 & ~n662 ;
  assign n664 = ~n647 & n662 ;
  assign n665 = ~n663 & ~n664 ;
  assign n666 = ~n626 & ~n665 ;
  assign n667 = ~n625 & ~n666 ;
  assign n668 = n617 & n667 ;
  assign n669 = ~n617 & ~n667 ;
  assign n670 = ~n645 & ~n663 ;
  assign n671 = ~n634 & ~n640 ;
  assign n672 = ~n670 & n671 ;
  assign n673 = n670 & ~n671 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~n655 & ~n661 ;
  assign n676 = n674 & n675 ;
  assign n677 = ~n674 & ~n675 ;
  assign n678 = ~n676 & ~n677 ;
  assign n679 = ~n669 & n678 ;
  assign n680 = ~n668 & ~n679 ;
  assign n681 = ~n615 & ~n680 ;
  assign n682 = n615 & n680 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = ~n672 & ~n676 ;
  assign n685 = n683 & ~n684 ;
  assign n686 = ~n681 & ~n685 ;
  assign n687 = ~n683 & n684 ;
  assign n688 = ~n685 & ~n687 ;
  assign n689 = ~x225 & ~x257 ;
  assign n690 = x225 & x257 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = ~n625 & ~n626 ;
  assign n693 = ~n665 & n692 ;
  assign n694 = n665 & ~n692 ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = ~n691 & ~n695 ;
  assign n697 = n691 & n695 ;
  assign n698 = ~x232 & ~x264 ;
  assign n699 = x232 & x264 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~x231 & ~x263 ;
  assign n702 = x231 & x263 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~n700 & ~n703 ;
  assign n705 = n700 & n703 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~x233 & ~x265 ;
  assign n708 = x233 & x265 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~n706 & ~n709 ;
  assign n711 = n706 & n709 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = ~x227 & ~x259 ;
  assign n714 = x227 & x259 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~n712 & ~n715 ;
  assign n717 = n712 & n715 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~x229 & ~x261 ;
  assign n720 = x229 & x261 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~x228 & ~x260 ;
  assign n723 = x228 & x260 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = ~n721 & ~n724 ;
  assign n726 = n721 & n724 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = ~x230 & ~x262 ;
  assign n729 = x230 & x262 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n727 & ~n730 ;
  assign n732 = n727 & n730 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = n718 & ~n733 ;
  assign n735 = ~n718 & n733 ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = ~x239 & ~x271 ;
  assign n738 = x239 & x271 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = ~x238 & ~x270 ;
  assign n741 = x238 & x270 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = ~n739 & ~n742 ;
  assign n744 = n739 & n742 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = ~x240 & ~x272 ;
  assign n747 = x240 & x272 ;
  assign n748 = ~n746 & ~n747 ;
  assign n749 = ~n745 & ~n748 ;
  assign n750 = n745 & n748 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~x234 & ~x266 ;
  assign n753 = x234 & x266 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~n751 & ~n754 ;
  assign n756 = n751 & n754 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = ~x236 & ~x268 ;
  assign n759 = x236 & x268 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = ~x235 & ~x267 ;
  assign n762 = x235 & x267 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~n760 & ~n763 ;
  assign n765 = n760 & n763 ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = ~x237 & ~x269 ;
  assign n768 = x237 & x269 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~n766 & ~n769 ;
  assign n771 = n766 & n769 ;
  assign n772 = ~n770 & ~n771 ;
  assign n773 = n757 & ~n772 ;
  assign n774 = ~n757 & n772 ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = ~x226 & ~x258 ;
  assign n777 = x226 & x258 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = n775 & ~n778 ;
  assign n780 = ~n775 & n778 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = n736 & n781 ;
  assign n783 = ~n736 & ~n781 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~n697 & n784 ;
  assign n786 = ~n696 & ~n785 ;
  assign n787 = ~n668 & ~n669 ;
  assign n788 = ~n678 & n787 ;
  assign n789 = n678 & ~n787 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = n786 & n790 ;
  assign n792 = ~n786 & ~n790 ;
  assign n793 = ~n716 & ~n734 ;
  assign n794 = ~n705 & ~n711 ;
  assign n795 = ~n793 & n794 ;
  assign n796 = n793 & ~n794 ;
  assign n797 = ~n795 & ~n796 ;
  assign n798 = ~n726 & ~n732 ;
  assign n799 = n797 & n798 ;
  assign n800 = ~n797 & ~n798 ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = ~n755 & ~n773 ;
  assign n803 = ~n744 & ~n750 ;
  assign n804 = ~n802 & n803 ;
  assign n805 = n802 & ~n803 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~n765 & ~n771 ;
  assign n808 = n806 & n807 ;
  assign n809 = ~n806 & ~n807 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n779 & ~n782 ;
  assign n812 = n810 & ~n811 ;
  assign n813 = ~n810 & n811 ;
  assign n814 = ~n812 & ~n813 ;
  assign n815 = n801 & n814 ;
  assign n816 = ~n801 & ~n814 ;
  assign n817 = ~n815 & ~n816 ;
  assign n818 = ~n792 & ~n817 ;
  assign n819 = ~n791 & ~n818 ;
  assign n820 = ~n688 & ~n819 ;
  assign n821 = n688 & n819 ;
  assign n822 = ~n801 & ~n812 ;
  assign n823 = ~n813 & ~n822 ;
  assign n824 = ~n804 & ~n808 ;
  assign n825 = n823 & ~n824 ;
  assign n826 = ~n823 & n824 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = ~n795 & ~n799 ;
  assign n829 = n827 & ~n828 ;
  assign n830 = ~n827 & n828 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = ~n821 & ~n831 ;
  assign n833 = ~n820 & ~n832 ;
  assign n834 = ~n686 & n833 ;
  assign n835 = n686 & ~n833 ;
  assign n836 = ~n834 & ~n835 ;
  assign n837 = ~n825 & ~n829 ;
  assign n838 = n836 & ~n837 ;
  assign n839 = ~n834 & ~n838 ;
  assign n840 = ~n836 & n837 ;
  assign n841 = ~n838 & ~n840 ;
  assign n842 = ~x224 & ~x256 ;
  assign n843 = x224 & x256 ;
  assign n844 = ~n842 & ~n843 ;
  assign n845 = ~n696 & ~n697 ;
  assign n846 = n784 & n845 ;
  assign n847 = ~n784 & ~n845 ;
  assign n848 = ~n846 & ~n847 ;
  assign n849 = n844 & ~n848 ;
  assign n850 = ~n791 & ~n792 ;
  assign n851 = ~n817 & n850 ;
  assign n852 = n817 & ~n850 ;
  assign n853 = ~n851 & ~n852 ;
  assign n854 = n849 & n853 ;
  assign n855 = ~n820 & ~n821 ;
  assign n856 = ~n831 & n855 ;
  assign n857 = n831 & ~n855 ;
  assign n858 = ~n856 & ~n857 ;
  assign n859 = n854 & n858 ;
  assign n860 = ~n841 & n859 ;
  assign n861 = n839 & n860 ;
  assign n862 = ~x222 & ~x286 ;
  assign n863 = x222 & x286 ;
  assign n864 = ~n862 & ~n863 ;
  assign n865 = ~x221 & ~x285 ;
  assign n866 = x221 & x285 ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = n864 & n867 ;
  assign n869 = ~n864 & ~n867 ;
  assign n870 = ~n868 & ~n869 ;
  assign n871 = ~x223 & ~x287 ;
  assign n872 = x223 & x287 ;
  assign n873 = ~n871 & ~n872 ;
  assign n874 = n870 & n873 ;
  assign n875 = ~n868 & ~n874 ;
  assign n876 = ~n870 & ~n873 ;
  assign n877 = ~n874 & ~n876 ;
  assign n878 = ~x217 & ~x281 ;
  assign n879 = x217 & x281 ;
  assign n880 = ~n878 & ~n879 ;
  assign n881 = n877 & n880 ;
  assign n882 = ~n877 & ~n880 ;
  assign n883 = ~x219 & ~x283 ;
  assign n884 = x219 & x283 ;
  assign n885 = ~n883 & ~n884 ;
  assign n886 = ~x218 & ~x282 ;
  assign n887 = x218 & x282 ;
  assign n888 = ~n886 & ~n887 ;
  assign n889 = ~n885 & ~n888 ;
  assign n890 = n885 & n888 ;
  assign n891 = ~n889 & ~n890 ;
  assign n892 = ~x220 & ~x284 ;
  assign n893 = x220 & x284 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = ~n891 & ~n894 ;
  assign n896 = n891 & n894 ;
  assign n897 = ~n895 & ~n896 ;
  assign n898 = ~n882 & n897 ;
  assign n899 = ~n881 & ~n898 ;
  assign n900 = n875 & n899 ;
  assign n901 = ~n875 & ~n899 ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = ~n890 & ~n896 ;
  assign n904 = n902 & n903 ;
  assign n905 = ~n900 & ~n904 ;
  assign n906 = ~n902 & ~n903 ;
  assign n907 = ~n904 & ~n906 ;
  assign n908 = ~n881 & ~n882 ;
  assign n909 = ~n897 & n908 ;
  assign n910 = n897 & ~n908 ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = ~x209 & ~x273 ;
  assign n913 = x209 & x273 ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = ~n911 & n914 ;
  assign n916 = n911 & ~n914 ;
  assign n917 = ~x215 & ~x279 ;
  assign n918 = x215 & x279 ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = ~x214 & ~x278 ;
  assign n921 = x214 & x278 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = ~n919 & ~n922 ;
  assign n924 = n919 & n922 ;
  assign n925 = ~n923 & ~n924 ;
  assign n926 = ~x216 & ~x280 ;
  assign n927 = x216 & x280 ;
  assign n928 = ~n926 & ~n927 ;
  assign n929 = ~n925 & ~n928 ;
  assign n930 = n925 & n928 ;
  assign n931 = ~n929 & ~n930 ;
  assign n932 = ~x210 & ~x274 ;
  assign n933 = x210 & x274 ;
  assign n934 = ~n932 & ~n933 ;
  assign n935 = ~n931 & ~n934 ;
  assign n936 = n931 & n934 ;
  assign n937 = ~n935 & ~n936 ;
  assign n938 = ~x212 & ~x276 ;
  assign n939 = x212 & x276 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = ~x211 & ~x275 ;
  assign n942 = x211 & x275 ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = ~n940 & ~n943 ;
  assign n945 = n940 & n943 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~x213 & ~x277 ;
  assign n948 = x213 & x277 ;
  assign n949 = ~n947 & ~n948 ;
  assign n950 = ~n946 & ~n949 ;
  assign n951 = n946 & n949 ;
  assign n952 = ~n950 & ~n951 ;
  assign n953 = n937 & ~n952 ;
  assign n954 = ~n937 & n952 ;
  assign n955 = ~n953 & ~n954 ;
  assign n956 = ~n916 & ~n955 ;
  assign n957 = ~n915 & ~n956 ;
  assign n958 = n907 & n957 ;
  assign n959 = ~n907 & ~n957 ;
  assign n960 = ~n935 & ~n953 ;
  assign n961 = ~n924 & ~n930 ;
  assign n962 = ~n960 & n961 ;
  assign n963 = n960 & ~n961 ;
  assign n964 = ~n962 & ~n963 ;
  assign n965 = ~n945 & ~n951 ;
  assign n966 = n964 & n965 ;
  assign n967 = ~n964 & ~n965 ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = ~n959 & n968 ;
  assign n970 = ~n958 & ~n969 ;
  assign n971 = ~n905 & ~n970 ;
  assign n972 = n905 & n970 ;
  assign n973 = ~n971 & ~n972 ;
  assign n974 = ~n962 & ~n966 ;
  assign n975 = n973 & ~n974 ;
  assign n976 = ~n971 & ~n975 ;
  assign n977 = ~n973 & n974 ;
  assign n978 = ~n975 & ~n977 ;
  assign n979 = ~x193 & ~x257 ;
  assign n980 = x193 & x257 ;
  assign n981 = ~n979 & ~n980 ;
  assign n982 = ~n915 & ~n916 ;
  assign n983 = ~n955 & n982 ;
  assign n984 = n955 & ~n982 ;
  assign n985 = ~n983 & ~n984 ;
  assign n986 = ~n981 & ~n985 ;
  assign n987 = n981 & n985 ;
  assign n988 = ~x200 & ~x264 ;
  assign n989 = x200 & x264 ;
  assign n990 = ~n988 & ~n989 ;
  assign n991 = ~x199 & ~x263 ;
  assign n992 = x199 & x263 ;
  assign n993 = ~n991 & ~n992 ;
  assign n994 = ~n990 & ~n993 ;
  assign n995 = n990 & n993 ;
  assign n996 = ~n994 & ~n995 ;
  assign n997 = ~x201 & ~x265 ;
  assign n998 = x201 & x265 ;
  assign n999 = ~n997 & ~n998 ;
  assign n1000 = ~n996 & ~n999 ;
  assign n1001 = n996 & n999 ;
  assign n1002 = ~n1000 & ~n1001 ;
  assign n1003 = ~x195 & ~x259 ;
  assign n1004 = x195 & x259 ;
  assign n1005 = ~n1003 & ~n1004 ;
  assign n1006 = ~n1002 & ~n1005 ;
  assign n1007 = n1002 & n1005 ;
  assign n1008 = ~n1006 & ~n1007 ;
  assign n1009 = ~x197 & ~x261 ;
  assign n1010 = x197 & x261 ;
  assign n1011 = ~n1009 & ~n1010 ;
  assign n1012 = ~x196 & ~x260 ;
  assign n1013 = x196 & x260 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = ~n1011 & ~n1014 ;
  assign n1016 = n1011 & n1014 ;
  assign n1017 = ~n1015 & ~n1016 ;
  assign n1018 = ~x198 & ~x262 ;
  assign n1019 = x198 & x262 ;
  assign n1020 = ~n1018 & ~n1019 ;
  assign n1021 = ~n1017 & ~n1020 ;
  assign n1022 = n1017 & n1020 ;
  assign n1023 = ~n1021 & ~n1022 ;
  assign n1024 = n1008 & ~n1023 ;
  assign n1025 = ~n1008 & n1023 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~x207 & ~x271 ;
  assign n1028 = x207 & x271 ;
  assign n1029 = ~n1027 & ~n1028 ;
  assign n1030 = ~x206 & ~x270 ;
  assign n1031 = x206 & x270 ;
  assign n1032 = ~n1030 & ~n1031 ;
  assign n1033 = ~n1029 & ~n1032 ;
  assign n1034 = n1029 & n1032 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1036 = ~x208 & ~x272 ;
  assign n1037 = x208 & x272 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = ~n1035 & ~n1038 ;
  assign n1040 = n1035 & n1038 ;
  assign n1041 = ~n1039 & ~n1040 ;
  assign n1042 = ~x202 & ~x266 ;
  assign n1043 = x202 & x266 ;
  assign n1044 = ~n1042 & ~n1043 ;
  assign n1045 = ~n1041 & ~n1044 ;
  assign n1046 = n1041 & n1044 ;
  assign n1047 = ~n1045 & ~n1046 ;
  assign n1048 = ~x204 & ~x268 ;
  assign n1049 = x204 & x268 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = ~x203 & ~x267 ;
  assign n1052 = x203 & x267 ;
  assign n1053 = ~n1051 & ~n1052 ;
  assign n1054 = ~n1050 & ~n1053 ;
  assign n1055 = n1050 & n1053 ;
  assign n1056 = ~n1054 & ~n1055 ;
  assign n1057 = ~x205 & ~x269 ;
  assign n1058 = x205 & x269 ;
  assign n1059 = ~n1057 & ~n1058 ;
  assign n1060 = ~n1056 & ~n1059 ;
  assign n1061 = n1056 & n1059 ;
  assign n1062 = ~n1060 & ~n1061 ;
  assign n1063 = n1047 & ~n1062 ;
  assign n1064 = ~n1047 & n1062 ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = ~x194 & ~x258 ;
  assign n1067 = x194 & x258 ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1069 = n1065 & ~n1068 ;
  assign n1070 = ~n1065 & n1068 ;
  assign n1071 = ~n1069 & ~n1070 ;
  assign n1072 = n1026 & n1071 ;
  assign n1073 = ~n1026 & ~n1071 ;
  assign n1074 = ~n1072 & ~n1073 ;
  assign n1075 = ~n987 & n1074 ;
  assign n1076 = ~n986 & ~n1075 ;
  assign n1077 = ~n958 & ~n959 ;
  assign n1078 = ~n968 & n1077 ;
  assign n1079 = n968 & ~n1077 ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1081 = n1076 & n1080 ;
  assign n1082 = ~n1076 & ~n1080 ;
  assign n1083 = ~n1006 & ~n1024 ;
  assign n1084 = ~n995 & ~n1001 ;
  assign n1085 = ~n1083 & n1084 ;
  assign n1086 = n1083 & ~n1084 ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1088 = ~n1016 & ~n1022 ;
  assign n1089 = n1087 & n1088 ;
  assign n1090 = ~n1087 & ~n1088 ;
  assign n1091 = ~n1089 & ~n1090 ;
  assign n1092 = ~n1045 & ~n1063 ;
  assign n1093 = ~n1034 & ~n1040 ;
  assign n1094 = ~n1092 & n1093 ;
  assign n1095 = n1092 & ~n1093 ;
  assign n1096 = ~n1094 & ~n1095 ;
  assign n1097 = ~n1055 & ~n1061 ;
  assign n1098 = n1096 & n1097 ;
  assign n1099 = ~n1096 & ~n1097 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = ~n1069 & ~n1072 ;
  assign n1102 = n1100 & ~n1101 ;
  assign n1103 = ~n1100 & n1101 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1105 = n1091 & n1104 ;
  assign n1106 = ~n1091 & ~n1104 ;
  assign n1107 = ~n1105 & ~n1106 ;
  assign n1108 = ~n1082 & ~n1107 ;
  assign n1109 = ~n1081 & ~n1108 ;
  assign n1110 = ~n978 & ~n1109 ;
  assign n1111 = n978 & n1109 ;
  assign n1112 = ~n1091 & ~n1102 ;
  assign n1113 = ~n1103 & ~n1112 ;
  assign n1114 = ~n1094 & ~n1098 ;
  assign n1115 = n1113 & ~n1114 ;
  assign n1116 = ~n1113 & n1114 ;
  assign n1117 = ~n1115 & ~n1116 ;
  assign n1118 = ~n1085 & ~n1089 ;
  assign n1119 = n1117 & ~n1118 ;
  assign n1120 = ~n1117 & n1118 ;
  assign n1121 = ~n1119 & ~n1120 ;
  assign n1122 = ~n1111 & ~n1121 ;
  assign n1123 = ~n1110 & ~n1122 ;
  assign n1124 = ~n976 & n1123 ;
  assign n1125 = n976 & ~n1123 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = ~n1115 & ~n1119 ;
  assign n1128 = n1126 & ~n1127 ;
  assign n1129 = ~n1124 & ~n1128 ;
  assign n1130 = ~n1126 & n1127 ;
  assign n1131 = ~n1128 & ~n1130 ;
  assign n1132 = ~x192 & ~x256 ;
  assign n1133 = x192 & x256 ;
  assign n1134 = ~n1132 & ~n1133 ;
  assign n1135 = ~n986 & ~n987 ;
  assign n1136 = n1074 & n1135 ;
  assign n1137 = ~n1074 & ~n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = n1134 & ~n1138 ;
  assign n1140 = ~n1081 & ~n1082 ;
  assign n1141 = ~n1107 & n1140 ;
  assign n1142 = n1107 & ~n1140 ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = n1139 & n1143 ;
  assign n1145 = ~n1110 & ~n1111 ;
  assign n1146 = ~n1121 & n1145 ;
  assign n1147 = n1121 & ~n1145 ;
  assign n1148 = ~n1146 & ~n1147 ;
  assign n1149 = n1144 & n1148 ;
  assign n1150 = ~n1131 & n1149 ;
  assign n1151 = n1129 & n1150 ;
  assign n1152 = ~n861 & ~n1151 ;
  assign n1153 = ~x190 & ~x286 ;
  assign n1154 = x190 & x286 ;
  assign n1155 = ~n1153 & ~n1154 ;
  assign n1156 = ~x189 & ~x285 ;
  assign n1157 = x189 & x285 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1159 = n1155 & n1158 ;
  assign n1160 = ~n1155 & ~n1158 ;
  assign n1161 = ~n1159 & ~n1160 ;
  assign n1162 = ~x191 & ~x287 ;
  assign n1163 = x191 & x287 ;
  assign n1164 = ~n1162 & ~n1163 ;
  assign n1165 = ~n1161 & ~n1164 ;
  assign n1166 = n1161 & n1164 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = ~x185 & ~x281 ;
  assign n1169 = x185 & x281 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = ~n1167 & ~n1170 ;
  assign n1172 = n1167 & n1170 ;
  assign n1173 = ~n1171 & ~n1172 ;
  assign n1174 = ~x187 & ~x283 ;
  assign n1175 = x187 & x283 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1177 = ~x186 & ~x282 ;
  assign n1178 = x186 & x282 ;
  assign n1179 = ~n1177 & ~n1178 ;
  assign n1180 = ~n1176 & ~n1179 ;
  assign n1181 = n1176 & n1179 ;
  assign n1182 = ~n1180 & ~n1181 ;
  assign n1183 = ~x188 & ~x284 ;
  assign n1184 = x188 & x284 ;
  assign n1185 = ~n1183 & ~n1184 ;
  assign n1186 = ~n1182 & ~n1185 ;
  assign n1187 = n1182 & n1185 ;
  assign n1188 = ~n1186 & ~n1187 ;
  assign n1189 = n1173 & ~n1188 ;
  assign n1190 = ~n1171 & ~n1189 ;
  assign n1191 = ~n1159 & ~n1166 ;
  assign n1192 = ~n1190 & n1191 ;
  assign n1193 = n1190 & ~n1191 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = ~n1181 & ~n1187 ;
  assign n1196 = n1194 & n1195 ;
  assign n1197 = ~n1192 & ~n1196 ;
  assign n1198 = ~n1194 & ~n1195 ;
  assign n1199 = ~n1196 & ~n1198 ;
  assign n1200 = ~n1173 & n1188 ;
  assign n1201 = ~n1189 & ~n1200 ;
  assign n1202 = ~x177 & ~x273 ;
  assign n1203 = x177 & x273 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1205 = n1201 & ~n1204 ;
  assign n1206 = ~x183 & ~x279 ;
  assign n1207 = x183 & x279 ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1209 = ~x182 & ~x278 ;
  assign n1210 = x182 & x278 ;
  assign n1211 = ~n1209 & ~n1210 ;
  assign n1212 = ~n1208 & ~n1211 ;
  assign n1213 = n1208 & n1211 ;
  assign n1214 = ~n1212 & ~n1213 ;
  assign n1215 = ~x184 & ~x280 ;
  assign n1216 = x184 & x280 ;
  assign n1217 = ~n1215 & ~n1216 ;
  assign n1218 = ~n1214 & ~n1217 ;
  assign n1219 = n1214 & n1217 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = ~x178 & ~x274 ;
  assign n1222 = x178 & x274 ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = ~n1220 & ~n1223 ;
  assign n1225 = n1220 & n1223 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1227 = ~x180 & ~x276 ;
  assign n1228 = x180 & x276 ;
  assign n1229 = ~n1227 & ~n1228 ;
  assign n1230 = ~x179 & ~x275 ;
  assign n1231 = x179 & x275 ;
  assign n1232 = ~n1230 & ~n1231 ;
  assign n1233 = ~n1229 & ~n1232 ;
  assign n1234 = n1229 & n1232 ;
  assign n1235 = ~n1233 & ~n1234 ;
  assign n1236 = ~x181 & ~x277 ;
  assign n1237 = x181 & x277 ;
  assign n1238 = ~n1236 & ~n1237 ;
  assign n1239 = ~n1235 & ~n1238 ;
  assign n1240 = n1235 & n1238 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = n1226 & ~n1241 ;
  assign n1243 = ~n1226 & n1241 ;
  assign n1244 = ~n1242 & ~n1243 ;
  assign n1245 = ~n1201 & n1204 ;
  assign n1246 = ~n1205 & ~n1245 ;
  assign n1247 = n1244 & n1246 ;
  assign n1248 = ~n1205 & ~n1247 ;
  assign n1249 = n1199 & ~n1248 ;
  assign n1250 = ~n1224 & ~n1242 ;
  assign n1251 = ~n1213 & ~n1219 ;
  assign n1252 = ~n1250 & n1251 ;
  assign n1253 = n1250 & ~n1251 ;
  assign n1254 = ~n1252 & ~n1253 ;
  assign n1255 = ~n1234 & ~n1240 ;
  assign n1256 = n1254 & n1255 ;
  assign n1257 = ~n1254 & ~n1255 ;
  assign n1258 = ~n1256 & ~n1257 ;
  assign n1259 = ~n1199 & n1248 ;
  assign n1260 = ~n1249 & ~n1259 ;
  assign n1261 = n1258 & n1260 ;
  assign n1262 = ~n1249 & ~n1261 ;
  assign n1263 = ~n1197 & ~n1262 ;
  assign n1264 = n1197 & n1262 ;
  assign n1265 = ~n1263 & ~n1264 ;
  assign n1266 = ~n1252 & ~n1256 ;
  assign n1267 = n1265 & ~n1266 ;
  assign n1268 = ~n1263 & ~n1267 ;
  assign n1269 = ~n1265 & n1266 ;
  assign n1270 = ~n1267 & ~n1269 ;
  assign n1271 = ~n1258 & ~n1260 ;
  assign n1272 = ~n1261 & ~n1271 ;
  assign n1273 = ~n1244 & ~n1246 ;
  assign n1274 = ~n1247 & ~n1273 ;
  assign n1275 = ~x161 & ~x257 ;
  assign n1276 = x161 & x257 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = n1274 & ~n1277 ;
  assign n1279 = ~x168 & ~x264 ;
  assign n1280 = x168 & x264 ;
  assign n1281 = ~n1279 & ~n1280 ;
  assign n1282 = ~x167 & ~x263 ;
  assign n1283 = x167 & x263 ;
  assign n1284 = ~n1282 & ~n1283 ;
  assign n1285 = ~n1281 & ~n1284 ;
  assign n1286 = n1281 & n1284 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = ~x169 & ~x265 ;
  assign n1289 = x169 & x265 ;
  assign n1290 = ~n1288 & ~n1289 ;
  assign n1291 = ~n1287 & ~n1290 ;
  assign n1292 = n1287 & n1290 ;
  assign n1293 = ~n1291 & ~n1292 ;
  assign n1294 = ~x163 & ~x259 ;
  assign n1295 = x163 & x259 ;
  assign n1296 = ~n1294 & ~n1295 ;
  assign n1297 = ~n1293 & ~n1296 ;
  assign n1298 = n1293 & n1296 ;
  assign n1299 = ~n1297 & ~n1298 ;
  assign n1300 = ~x165 & ~x261 ;
  assign n1301 = x165 & x261 ;
  assign n1302 = ~n1300 & ~n1301 ;
  assign n1303 = ~x164 & ~x260 ;
  assign n1304 = x164 & x260 ;
  assign n1305 = ~n1303 & ~n1304 ;
  assign n1306 = ~n1302 & ~n1305 ;
  assign n1307 = n1302 & n1305 ;
  assign n1308 = ~n1306 & ~n1307 ;
  assign n1309 = ~x166 & ~x262 ;
  assign n1310 = x166 & x262 ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1312 = ~n1308 & ~n1311 ;
  assign n1313 = n1308 & n1311 ;
  assign n1314 = ~n1312 & ~n1313 ;
  assign n1315 = n1299 & ~n1314 ;
  assign n1316 = ~n1299 & n1314 ;
  assign n1317 = ~n1315 & ~n1316 ;
  assign n1318 = ~x175 & ~x271 ;
  assign n1319 = x175 & x271 ;
  assign n1320 = ~n1318 & ~n1319 ;
  assign n1321 = ~x174 & ~x270 ;
  assign n1322 = x174 & x270 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = ~n1320 & ~n1323 ;
  assign n1325 = n1320 & n1323 ;
  assign n1326 = ~n1324 & ~n1325 ;
  assign n1327 = ~x176 & ~x272 ;
  assign n1328 = x176 & x272 ;
  assign n1329 = ~n1327 & ~n1328 ;
  assign n1330 = ~n1326 & ~n1329 ;
  assign n1331 = n1326 & n1329 ;
  assign n1332 = ~n1330 & ~n1331 ;
  assign n1333 = ~x170 & ~x266 ;
  assign n1334 = x170 & x266 ;
  assign n1335 = ~n1333 & ~n1334 ;
  assign n1336 = ~n1332 & ~n1335 ;
  assign n1337 = n1332 & n1335 ;
  assign n1338 = ~n1336 & ~n1337 ;
  assign n1339 = ~x172 & ~x268 ;
  assign n1340 = x172 & x268 ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1342 = ~x171 & ~x267 ;
  assign n1343 = x171 & x267 ;
  assign n1344 = ~n1342 & ~n1343 ;
  assign n1345 = ~n1341 & ~n1344 ;
  assign n1346 = n1341 & n1344 ;
  assign n1347 = ~n1345 & ~n1346 ;
  assign n1348 = ~x173 & ~x269 ;
  assign n1349 = x173 & x269 ;
  assign n1350 = ~n1348 & ~n1349 ;
  assign n1351 = ~n1347 & ~n1350 ;
  assign n1352 = n1347 & n1350 ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = n1338 & ~n1353 ;
  assign n1355 = ~n1338 & n1353 ;
  assign n1356 = ~n1354 & ~n1355 ;
  assign n1357 = ~x162 & ~x258 ;
  assign n1358 = x162 & x258 ;
  assign n1359 = ~n1357 & ~n1358 ;
  assign n1360 = n1356 & ~n1359 ;
  assign n1361 = ~n1356 & n1359 ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = n1317 & n1362 ;
  assign n1364 = ~n1317 & ~n1362 ;
  assign n1365 = ~n1363 & ~n1364 ;
  assign n1366 = ~n1274 & n1277 ;
  assign n1367 = ~n1278 & ~n1366 ;
  assign n1368 = n1365 & n1367 ;
  assign n1369 = ~n1278 & ~n1368 ;
  assign n1370 = n1272 & ~n1369 ;
  assign n1371 = ~n1297 & ~n1315 ;
  assign n1372 = ~n1286 & ~n1292 ;
  assign n1373 = ~n1371 & n1372 ;
  assign n1374 = n1371 & ~n1372 ;
  assign n1375 = ~n1373 & ~n1374 ;
  assign n1376 = ~n1307 & ~n1313 ;
  assign n1377 = n1375 & n1376 ;
  assign n1378 = ~n1375 & ~n1376 ;
  assign n1379 = ~n1377 & ~n1378 ;
  assign n1380 = ~n1336 & ~n1354 ;
  assign n1381 = ~n1325 & ~n1331 ;
  assign n1382 = ~n1380 & n1381 ;
  assign n1383 = n1380 & ~n1381 ;
  assign n1384 = ~n1382 & ~n1383 ;
  assign n1385 = ~n1346 & ~n1352 ;
  assign n1386 = n1384 & n1385 ;
  assign n1387 = ~n1384 & ~n1385 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = ~n1360 & ~n1363 ;
  assign n1390 = n1388 & ~n1389 ;
  assign n1391 = ~n1388 & n1389 ;
  assign n1392 = ~n1390 & ~n1391 ;
  assign n1393 = n1379 & n1392 ;
  assign n1394 = ~n1379 & ~n1392 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = ~n1272 & n1369 ;
  assign n1397 = ~n1370 & ~n1396 ;
  assign n1398 = n1395 & n1397 ;
  assign n1399 = ~n1370 & ~n1398 ;
  assign n1400 = n1270 & ~n1399 ;
  assign n1401 = ~n1382 & ~n1386 ;
  assign n1402 = ~n1390 & ~n1393 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = n1401 & n1402 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~n1373 & ~n1377 ;
  assign n1407 = n1405 & ~n1406 ;
  assign n1408 = ~n1405 & n1406 ;
  assign n1409 = ~n1407 & ~n1408 ;
  assign n1410 = ~n1270 & n1399 ;
  assign n1411 = ~n1400 & ~n1410 ;
  assign n1412 = n1409 & n1411 ;
  assign n1413 = ~n1400 & ~n1412 ;
  assign n1414 = ~n1268 & ~n1413 ;
  assign n1415 = n1268 & n1413 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~n1403 & ~n1407 ;
  assign n1418 = n1416 & ~n1417 ;
  assign n1419 = ~n1414 & ~n1418 ;
  assign n1420 = ~n1416 & n1417 ;
  assign n1421 = ~n1418 & ~n1420 ;
  assign n1422 = ~n1409 & ~n1411 ;
  assign n1423 = ~n1412 & ~n1422 ;
  assign n1424 = ~n1395 & ~n1397 ;
  assign n1425 = ~n1398 & ~n1424 ;
  assign n1426 = ~n1365 & ~n1367 ;
  assign n1427 = ~n1368 & ~n1426 ;
  assign n1428 = ~x160 & ~x256 ;
  assign n1429 = x160 & x256 ;
  assign n1430 = ~n1428 & ~n1429 ;
  assign n1431 = ~n1427 & n1430 ;
  assign n1432 = ~n1425 & n1431 ;
  assign n1433 = ~n1423 & n1432 ;
  assign n1434 = ~n1421 & n1433 ;
  assign n1435 = n1419 & n1434 ;
  assign n1436 = ~n1152 & n1435 ;
  assign n1437 = n861 & n1151 ;
  assign n1438 = ~n1435 & n1437 ;
  assign n1439 = ~n1436 & ~n1438 ;
  assign n1440 = n1152 & ~n1435 ;
  assign n1441 = ~x158 & ~x286 ;
  assign n1442 = x158 & x286 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = ~x157 & ~x285 ;
  assign n1445 = x157 & x285 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = n1443 & n1446 ;
  assign n1448 = ~n1443 & ~n1446 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1450 = ~x159 & ~x287 ;
  assign n1451 = x159 & x287 ;
  assign n1452 = ~n1450 & ~n1451 ;
  assign n1453 = ~n1449 & ~n1452 ;
  assign n1454 = n1449 & n1452 ;
  assign n1455 = ~n1453 & ~n1454 ;
  assign n1456 = ~x153 & ~x281 ;
  assign n1457 = x153 & x281 ;
  assign n1458 = ~n1456 & ~n1457 ;
  assign n1459 = ~n1455 & ~n1458 ;
  assign n1460 = n1455 & n1458 ;
  assign n1461 = ~n1459 & ~n1460 ;
  assign n1462 = ~x155 & ~x283 ;
  assign n1463 = x155 & x283 ;
  assign n1464 = ~n1462 & ~n1463 ;
  assign n1465 = ~x154 & ~x282 ;
  assign n1466 = x154 & x282 ;
  assign n1467 = ~n1465 & ~n1466 ;
  assign n1468 = ~n1464 & ~n1467 ;
  assign n1469 = n1464 & n1467 ;
  assign n1470 = ~n1468 & ~n1469 ;
  assign n1471 = ~x156 & ~x284 ;
  assign n1472 = x156 & x284 ;
  assign n1473 = ~n1471 & ~n1472 ;
  assign n1474 = ~n1470 & ~n1473 ;
  assign n1475 = n1470 & n1473 ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = n1461 & ~n1476 ;
  assign n1478 = ~n1459 & ~n1477 ;
  assign n1479 = ~n1447 & ~n1454 ;
  assign n1480 = ~n1478 & n1479 ;
  assign n1481 = n1478 & ~n1479 ;
  assign n1482 = ~n1480 & ~n1481 ;
  assign n1483 = ~n1469 & ~n1475 ;
  assign n1484 = n1482 & n1483 ;
  assign n1485 = ~n1480 & ~n1484 ;
  assign n1486 = ~n1482 & ~n1483 ;
  assign n1487 = ~n1484 & ~n1486 ;
  assign n1488 = ~n1461 & n1476 ;
  assign n1489 = ~n1477 & ~n1488 ;
  assign n1490 = ~x145 & ~x273 ;
  assign n1491 = x145 & x273 ;
  assign n1492 = ~n1490 & ~n1491 ;
  assign n1493 = n1489 & ~n1492 ;
  assign n1494 = ~x151 & ~x279 ;
  assign n1495 = x151 & x279 ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = ~x150 & ~x278 ;
  assign n1498 = x150 & x278 ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = ~n1496 & ~n1499 ;
  assign n1501 = n1496 & n1499 ;
  assign n1502 = ~n1500 & ~n1501 ;
  assign n1503 = ~x152 & ~x280 ;
  assign n1504 = x152 & x280 ;
  assign n1505 = ~n1503 & ~n1504 ;
  assign n1506 = ~n1502 & ~n1505 ;
  assign n1507 = n1502 & n1505 ;
  assign n1508 = ~n1506 & ~n1507 ;
  assign n1509 = ~x146 & ~x274 ;
  assign n1510 = x146 & x274 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = ~n1508 & ~n1511 ;
  assign n1513 = n1508 & n1511 ;
  assign n1514 = ~n1512 & ~n1513 ;
  assign n1515 = ~x148 & ~x276 ;
  assign n1516 = x148 & x276 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = ~x147 & ~x275 ;
  assign n1519 = x147 & x275 ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = ~n1517 & ~n1520 ;
  assign n1522 = n1517 & n1520 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = ~x149 & ~x277 ;
  assign n1525 = x149 & x277 ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = ~n1523 & ~n1526 ;
  assign n1528 = n1523 & n1526 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1530 = n1514 & ~n1529 ;
  assign n1531 = ~n1514 & n1529 ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1533 = ~n1489 & n1492 ;
  assign n1534 = ~n1493 & ~n1533 ;
  assign n1535 = n1532 & n1534 ;
  assign n1536 = ~n1493 & ~n1535 ;
  assign n1537 = n1487 & ~n1536 ;
  assign n1538 = ~n1512 & ~n1530 ;
  assign n1539 = ~n1501 & ~n1507 ;
  assign n1540 = ~n1538 & n1539 ;
  assign n1541 = n1538 & ~n1539 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = ~n1522 & ~n1528 ;
  assign n1544 = n1542 & n1543 ;
  assign n1545 = ~n1542 & ~n1543 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = ~n1487 & n1536 ;
  assign n1548 = ~n1537 & ~n1547 ;
  assign n1549 = n1546 & n1548 ;
  assign n1550 = ~n1537 & ~n1549 ;
  assign n1551 = ~n1485 & ~n1550 ;
  assign n1552 = n1485 & n1550 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = ~n1540 & ~n1544 ;
  assign n1555 = n1553 & ~n1554 ;
  assign n1556 = ~n1551 & ~n1555 ;
  assign n1557 = ~n1553 & n1554 ;
  assign n1558 = ~n1555 & ~n1557 ;
  assign n1559 = ~n1546 & ~n1548 ;
  assign n1560 = ~n1549 & ~n1559 ;
  assign n1561 = ~n1532 & ~n1534 ;
  assign n1562 = ~n1535 & ~n1561 ;
  assign n1563 = ~x129 & ~x257 ;
  assign n1564 = x129 & x257 ;
  assign n1565 = ~n1563 & ~n1564 ;
  assign n1566 = n1562 & ~n1565 ;
  assign n1567 = ~x136 & ~x264 ;
  assign n1568 = x136 & x264 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = ~x135 & ~x263 ;
  assign n1571 = x135 & x263 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = ~n1569 & ~n1572 ;
  assign n1574 = n1569 & n1572 ;
  assign n1575 = ~n1573 & ~n1574 ;
  assign n1576 = ~x137 & ~x265 ;
  assign n1577 = x137 & x265 ;
  assign n1578 = ~n1576 & ~n1577 ;
  assign n1579 = ~n1575 & ~n1578 ;
  assign n1580 = n1575 & n1578 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = ~x131 & ~x259 ;
  assign n1583 = x131 & x259 ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1585 = ~n1581 & ~n1584 ;
  assign n1586 = n1581 & n1584 ;
  assign n1587 = ~n1585 & ~n1586 ;
  assign n1588 = ~x133 & ~x261 ;
  assign n1589 = x133 & x261 ;
  assign n1590 = ~n1588 & ~n1589 ;
  assign n1591 = ~x132 & ~x260 ;
  assign n1592 = x132 & x260 ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = ~n1590 & ~n1593 ;
  assign n1595 = n1590 & n1593 ;
  assign n1596 = ~n1594 & ~n1595 ;
  assign n1597 = ~x134 & ~x262 ;
  assign n1598 = x134 & x262 ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = ~n1596 & ~n1599 ;
  assign n1601 = n1596 & n1599 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = n1587 & ~n1602 ;
  assign n1604 = ~n1587 & n1602 ;
  assign n1605 = ~n1603 & ~n1604 ;
  assign n1606 = ~x143 & ~x271 ;
  assign n1607 = x143 & x271 ;
  assign n1608 = ~n1606 & ~n1607 ;
  assign n1609 = ~x142 & ~x270 ;
  assign n1610 = x142 & x270 ;
  assign n1611 = ~n1609 & ~n1610 ;
  assign n1612 = ~n1608 & ~n1611 ;
  assign n1613 = n1608 & n1611 ;
  assign n1614 = ~n1612 & ~n1613 ;
  assign n1615 = ~x144 & ~x272 ;
  assign n1616 = x144 & x272 ;
  assign n1617 = ~n1615 & ~n1616 ;
  assign n1618 = ~n1614 & ~n1617 ;
  assign n1619 = n1614 & n1617 ;
  assign n1620 = ~n1618 & ~n1619 ;
  assign n1621 = ~x138 & ~x266 ;
  assign n1622 = x138 & x266 ;
  assign n1623 = ~n1621 & ~n1622 ;
  assign n1624 = ~n1620 & ~n1623 ;
  assign n1625 = n1620 & n1623 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1627 = ~x140 & ~x268 ;
  assign n1628 = x140 & x268 ;
  assign n1629 = ~n1627 & ~n1628 ;
  assign n1630 = ~x139 & ~x267 ;
  assign n1631 = x139 & x267 ;
  assign n1632 = ~n1630 & ~n1631 ;
  assign n1633 = ~n1629 & ~n1632 ;
  assign n1634 = n1629 & n1632 ;
  assign n1635 = ~n1633 & ~n1634 ;
  assign n1636 = ~x141 & ~x269 ;
  assign n1637 = x141 & x269 ;
  assign n1638 = ~n1636 & ~n1637 ;
  assign n1639 = ~n1635 & ~n1638 ;
  assign n1640 = n1635 & n1638 ;
  assign n1641 = ~n1639 & ~n1640 ;
  assign n1642 = n1626 & ~n1641 ;
  assign n1643 = ~n1626 & n1641 ;
  assign n1644 = ~n1642 & ~n1643 ;
  assign n1645 = ~x130 & ~x258 ;
  assign n1646 = x130 & x258 ;
  assign n1647 = ~n1645 & ~n1646 ;
  assign n1648 = n1644 & ~n1647 ;
  assign n1649 = ~n1644 & n1647 ;
  assign n1650 = ~n1648 & ~n1649 ;
  assign n1651 = n1605 & n1650 ;
  assign n1652 = ~n1605 & ~n1650 ;
  assign n1653 = ~n1651 & ~n1652 ;
  assign n1654 = ~n1562 & n1565 ;
  assign n1655 = ~n1566 & ~n1654 ;
  assign n1656 = n1653 & n1655 ;
  assign n1657 = ~n1566 & ~n1656 ;
  assign n1658 = n1560 & ~n1657 ;
  assign n1659 = ~n1585 & ~n1603 ;
  assign n1660 = ~n1574 & ~n1580 ;
  assign n1661 = ~n1659 & n1660 ;
  assign n1662 = n1659 & ~n1660 ;
  assign n1663 = ~n1661 & ~n1662 ;
  assign n1664 = ~n1595 & ~n1601 ;
  assign n1665 = n1663 & n1664 ;
  assign n1666 = ~n1663 & ~n1664 ;
  assign n1667 = ~n1665 & ~n1666 ;
  assign n1668 = ~n1624 & ~n1642 ;
  assign n1669 = ~n1613 & ~n1619 ;
  assign n1670 = ~n1668 & n1669 ;
  assign n1671 = n1668 & ~n1669 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = ~n1634 & ~n1640 ;
  assign n1674 = n1672 & n1673 ;
  assign n1675 = ~n1672 & ~n1673 ;
  assign n1676 = ~n1674 & ~n1675 ;
  assign n1677 = ~n1648 & ~n1651 ;
  assign n1678 = n1676 & ~n1677 ;
  assign n1679 = ~n1676 & n1677 ;
  assign n1680 = ~n1678 & ~n1679 ;
  assign n1681 = n1667 & n1680 ;
  assign n1682 = ~n1667 & ~n1680 ;
  assign n1683 = ~n1681 & ~n1682 ;
  assign n1684 = ~n1560 & n1657 ;
  assign n1685 = ~n1658 & ~n1684 ;
  assign n1686 = n1683 & n1685 ;
  assign n1687 = ~n1658 & ~n1686 ;
  assign n1688 = n1558 & ~n1687 ;
  assign n1689 = ~n1670 & ~n1674 ;
  assign n1690 = ~n1678 & ~n1681 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = n1689 & n1690 ;
  assign n1693 = ~n1691 & ~n1692 ;
  assign n1694 = ~n1661 & ~n1665 ;
  assign n1695 = n1693 & ~n1694 ;
  assign n1696 = ~n1693 & n1694 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1698 = ~n1558 & n1687 ;
  assign n1699 = ~n1688 & ~n1698 ;
  assign n1700 = n1697 & n1699 ;
  assign n1701 = ~n1688 & ~n1700 ;
  assign n1702 = ~n1556 & ~n1701 ;
  assign n1703 = n1556 & n1701 ;
  assign n1704 = ~n1702 & ~n1703 ;
  assign n1705 = ~n1691 & ~n1695 ;
  assign n1706 = n1704 & ~n1705 ;
  assign n1707 = ~n1702 & ~n1706 ;
  assign n1708 = ~n1704 & n1705 ;
  assign n1709 = ~n1706 & ~n1708 ;
  assign n1710 = ~n1697 & ~n1699 ;
  assign n1711 = ~n1700 & ~n1710 ;
  assign n1712 = ~n1683 & ~n1685 ;
  assign n1713 = ~n1686 & ~n1712 ;
  assign n1714 = ~n1653 & ~n1655 ;
  assign n1715 = ~n1656 & ~n1714 ;
  assign n1716 = ~x128 & ~x256 ;
  assign n1717 = x128 & x256 ;
  assign n1718 = ~n1716 & ~n1717 ;
  assign n1719 = ~n1715 & n1718 ;
  assign n1720 = ~n1713 & n1719 ;
  assign n1721 = ~n1711 & n1720 ;
  assign n1722 = ~n1709 & n1721 ;
  assign n1723 = n1707 & n1722 ;
  assign n1724 = ~n1440 & n1723 ;
  assign n1725 = ~n1439 & n1724 ;
  assign n1726 = n1435 & n1437 ;
  assign n1727 = ~n1723 & n1726 ;
  assign n1728 = ~n1725 & ~n1727 ;
  assign n1729 = n1439 & ~n1724 ;
  assign n1730 = ~x126 & ~x286 ;
  assign n1731 = x126 & x286 ;
  assign n1732 = ~n1730 & ~n1731 ;
  assign n1733 = ~x125 & ~x285 ;
  assign n1734 = x125 & x285 ;
  assign n1735 = ~n1733 & ~n1734 ;
  assign n1736 = n1732 & n1735 ;
  assign n1737 = ~n1732 & ~n1735 ;
  assign n1738 = ~n1736 & ~n1737 ;
  assign n1739 = ~x127 & ~x287 ;
  assign n1740 = x127 & x287 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1738 & ~n1741 ;
  assign n1743 = n1738 & n1741 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = ~x121 & ~x281 ;
  assign n1746 = x121 & x281 ;
  assign n1747 = ~n1745 & ~n1746 ;
  assign n1748 = ~n1744 & ~n1747 ;
  assign n1749 = n1744 & n1747 ;
  assign n1750 = ~n1748 & ~n1749 ;
  assign n1751 = ~x123 & ~x283 ;
  assign n1752 = x123 & x283 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1754 = ~x122 & ~x282 ;
  assign n1755 = x122 & x282 ;
  assign n1756 = ~n1754 & ~n1755 ;
  assign n1757 = ~n1753 & ~n1756 ;
  assign n1758 = n1753 & n1756 ;
  assign n1759 = ~n1757 & ~n1758 ;
  assign n1760 = ~x124 & ~x284 ;
  assign n1761 = x124 & x284 ;
  assign n1762 = ~n1760 & ~n1761 ;
  assign n1763 = ~n1759 & ~n1762 ;
  assign n1764 = n1759 & n1762 ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1766 = n1750 & ~n1765 ;
  assign n1767 = ~n1748 & ~n1766 ;
  assign n1768 = ~n1736 & ~n1743 ;
  assign n1769 = ~n1767 & n1768 ;
  assign n1770 = n1767 & ~n1768 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = ~n1758 & ~n1764 ;
  assign n1773 = n1771 & n1772 ;
  assign n1774 = ~n1769 & ~n1773 ;
  assign n1775 = ~n1771 & ~n1772 ;
  assign n1776 = ~n1773 & ~n1775 ;
  assign n1777 = ~n1750 & n1765 ;
  assign n1778 = ~n1766 & ~n1777 ;
  assign n1779 = ~x113 & ~x273 ;
  assign n1780 = x113 & x273 ;
  assign n1781 = ~n1779 & ~n1780 ;
  assign n1782 = n1778 & ~n1781 ;
  assign n1783 = ~x119 & ~x279 ;
  assign n1784 = x119 & x279 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = ~x118 & ~x278 ;
  assign n1787 = x118 & x278 ;
  assign n1788 = ~n1786 & ~n1787 ;
  assign n1789 = ~n1785 & ~n1788 ;
  assign n1790 = n1785 & n1788 ;
  assign n1791 = ~n1789 & ~n1790 ;
  assign n1792 = ~x120 & ~x280 ;
  assign n1793 = x120 & x280 ;
  assign n1794 = ~n1792 & ~n1793 ;
  assign n1795 = ~n1791 & ~n1794 ;
  assign n1796 = n1791 & n1794 ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1798 = ~x114 & ~x274 ;
  assign n1799 = x114 & x274 ;
  assign n1800 = ~n1798 & ~n1799 ;
  assign n1801 = ~n1797 & ~n1800 ;
  assign n1802 = n1797 & n1800 ;
  assign n1803 = ~n1801 & ~n1802 ;
  assign n1804 = ~x116 & ~x276 ;
  assign n1805 = x116 & x276 ;
  assign n1806 = ~n1804 & ~n1805 ;
  assign n1807 = ~x115 & ~x275 ;
  assign n1808 = x115 & x275 ;
  assign n1809 = ~n1807 & ~n1808 ;
  assign n1810 = ~n1806 & ~n1809 ;
  assign n1811 = n1806 & n1809 ;
  assign n1812 = ~n1810 & ~n1811 ;
  assign n1813 = ~x117 & ~x277 ;
  assign n1814 = x117 & x277 ;
  assign n1815 = ~n1813 & ~n1814 ;
  assign n1816 = ~n1812 & ~n1815 ;
  assign n1817 = n1812 & n1815 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = n1803 & ~n1818 ;
  assign n1820 = ~n1803 & n1818 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1822 = ~n1778 & n1781 ;
  assign n1823 = ~n1782 & ~n1822 ;
  assign n1824 = n1821 & n1823 ;
  assign n1825 = ~n1782 & ~n1824 ;
  assign n1826 = n1776 & ~n1825 ;
  assign n1827 = ~n1801 & ~n1819 ;
  assign n1828 = ~n1790 & ~n1796 ;
  assign n1829 = ~n1827 & n1828 ;
  assign n1830 = n1827 & ~n1828 ;
  assign n1831 = ~n1829 & ~n1830 ;
  assign n1832 = ~n1811 & ~n1817 ;
  assign n1833 = n1831 & n1832 ;
  assign n1834 = ~n1831 & ~n1832 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = ~n1776 & n1825 ;
  assign n1837 = ~n1826 & ~n1836 ;
  assign n1838 = n1835 & n1837 ;
  assign n1839 = ~n1826 & ~n1838 ;
  assign n1840 = ~n1774 & ~n1839 ;
  assign n1841 = n1774 & n1839 ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = ~n1829 & ~n1833 ;
  assign n1844 = n1842 & ~n1843 ;
  assign n1845 = ~n1840 & ~n1844 ;
  assign n1846 = ~n1842 & n1843 ;
  assign n1847 = ~n1844 & ~n1846 ;
  assign n1848 = ~n1835 & ~n1837 ;
  assign n1849 = ~n1838 & ~n1848 ;
  assign n1850 = ~n1821 & ~n1823 ;
  assign n1851 = ~n1824 & ~n1850 ;
  assign n1852 = ~x97 & ~x257 ;
  assign n1853 = x97 & x257 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = n1851 & ~n1854 ;
  assign n1856 = ~x104 & ~x264 ;
  assign n1857 = x104 & x264 ;
  assign n1858 = ~n1856 & ~n1857 ;
  assign n1859 = ~x103 & ~x263 ;
  assign n1860 = x103 & x263 ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = ~n1858 & ~n1861 ;
  assign n1863 = n1858 & n1861 ;
  assign n1864 = ~n1862 & ~n1863 ;
  assign n1865 = ~x105 & ~x265 ;
  assign n1866 = x105 & x265 ;
  assign n1867 = ~n1865 & ~n1866 ;
  assign n1868 = ~n1864 & ~n1867 ;
  assign n1869 = n1864 & n1867 ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = ~x99 & ~x259 ;
  assign n1872 = x99 & x259 ;
  assign n1873 = ~n1871 & ~n1872 ;
  assign n1874 = ~n1870 & ~n1873 ;
  assign n1875 = n1870 & n1873 ;
  assign n1876 = ~n1874 & ~n1875 ;
  assign n1877 = ~x101 & ~x261 ;
  assign n1878 = x101 & x261 ;
  assign n1879 = ~n1877 & ~n1878 ;
  assign n1880 = ~x100 & ~x260 ;
  assign n1881 = x100 & x260 ;
  assign n1882 = ~n1880 & ~n1881 ;
  assign n1883 = ~n1879 & ~n1882 ;
  assign n1884 = n1879 & n1882 ;
  assign n1885 = ~n1883 & ~n1884 ;
  assign n1886 = ~x102 & ~x262 ;
  assign n1887 = x102 & x262 ;
  assign n1888 = ~n1886 & ~n1887 ;
  assign n1889 = ~n1885 & ~n1888 ;
  assign n1890 = n1885 & n1888 ;
  assign n1891 = ~n1889 & ~n1890 ;
  assign n1892 = n1876 & ~n1891 ;
  assign n1893 = ~n1876 & n1891 ;
  assign n1894 = ~n1892 & ~n1893 ;
  assign n1895 = ~x111 & ~x271 ;
  assign n1896 = x111 & x271 ;
  assign n1897 = ~n1895 & ~n1896 ;
  assign n1898 = ~x110 & ~x270 ;
  assign n1899 = x110 & x270 ;
  assign n1900 = ~n1898 & ~n1899 ;
  assign n1901 = ~n1897 & ~n1900 ;
  assign n1902 = n1897 & n1900 ;
  assign n1903 = ~n1901 & ~n1902 ;
  assign n1904 = ~x112 & ~x272 ;
  assign n1905 = x112 & x272 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1907 = ~n1903 & ~n1906 ;
  assign n1908 = n1903 & n1906 ;
  assign n1909 = ~n1907 & ~n1908 ;
  assign n1910 = ~x106 & ~x266 ;
  assign n1911 = x106 & x266 ;
  assign n1912 = ~n1910 & ~n1911 ;
  assign n1913 = ~n1909 & ~n1912 ;
  assign n1914 = n1909 & n1912 ;
  assign n1915 = ~n1913 & ~n1914 ;
  assign n1916 = ~x108 & ~x268 ;
  assign n1917 = x108 & x268 ;
  assign n1918 = ~n1916 & ~n1917 ;
  assign n1919 = ~x107 & ~x267 ;
  assign n1920 = x107 & x267 ;
  assign n1921 = ~n1919 & ~n1920 ;
  assign n1922 = ~n1918 & ~n1921 ;
  assign n1923 = n1918 & n1921 ;
  assign n1924 = ~n1922 & ~n1923 ;
  assign n1925 = ~x109 & ~x269 ;
  assign n1926 = x109 & x269 ;
  assign n1927 = ~n1925 & ~n1926 ;
  assign n1928 = ~n1924 & ~n1927 ;
  assign n1929 = n1924 & n1927 ;
  assign n1930 = ~n1928 & ~n1929 ;
  assign n1931 = n1915 & ~n1930 ;
  assign n1932 = ~n1915 & n1930 ;
  assign n1933 = ~n1931 & ~n1932 ;
  assign n1934 = ~x98 & ~x258 ;
  assign n1935 = x98 & x258 ;
  assign n1936 = ~n1934 & ~n1935 ;
  assign n1937 = n1933 & ~n1936 ;
  assign n1938 = ~n1933 & n1936 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = n1894 & n1939 ;
  assign n1941 = ~n1894 & ~n1939 ;
  assign n1942 = ~n1940 & ~n1941 ;
  assign n1943 = ~n1851 & n1854 ;
  assign n1944 = ~n1855 & ~n1943 ;
  assign n1945 = n1942 & n1944 ;
  assign n1946 = ~n1855 & ~n1945 ;
  assign n1947 = n1849 & ~n1946 ;
  assign n1948 = ~n1874 & ~n1892 ;
  assign n1949 = ~n1863 & ~n1869 ;
  assign n1950 = ~n1948 & n1949 ;
  assign n1951 = n1948 & ~n1949 ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1953 = ~n1884 & ~n1890 ;
  assign n1954 = n1952 & n1953 ;
  assign n1955 = ~n1952 & ~n1953 ;
  assign n1956 = ~n1954 & ~n1955 ;
  assign n1957 = ~n1913 & ~n1931 ;
  assign n1958 = ~n1902 & ~n1908 ;
  assign n1959 = ~n1957 & n1958 ;
  assign n1960 = n1957 & ~n1958 ;
  assign n1961 = ~n1959 & ~n1960 ;
  assign n1962 = ~n1923 & ~n1929 ;
  assign n1963 = n1961 & n1962 ;
  assign n1964 = ~n1961 & ~n1962 ;
  assign n1965 = ~n1963 & ~n1964 ;
  assign n1966 = ~n1937 & ~n1940 ;
  assign n1967 = n1965 & ~n1966 ;
  assign n1968 = ~n1965 & n1966 ;
  assign n1969 = ~n1967 & ~n1968 ;
  assign n1970 = n1956 & n1969 ;
  assign n1971 = ~n1956 & ~n1969 ;
  assign n1972 = ~n1970 & ~n1971 ;
  assign n1973 = ~n1849 & n1946 ;
  assign n1974 = ~n1947 & ~n1973 ;
  assign n1975 = n1972 & n1974 ;
  assign n1976 = ~n1947 & ~n1975 ;
  assign n1977 = n1847 & ~n1976 ;
  assign n1978 = ~n1959 & ~n1963 ;
  assign n1979 = ~n1967 & ~n1970 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = n1978 & n1979 ;
  assign n1982 = ~n1980 & ~n1981 ;
  assign n1983 = ~n1950 & ~n1954 ;
  assign n1984 = n1982 & ~n1983 ;
  assign n1985 = ~n1982 & n1983 ;
  assign n1986 = ~n1984 & ~n1985 ;
  assign n1987 = ~n1847 & n1976 ;
  assign n1988 = ~n1977 & ~n1987 ;
  assign n1989 = n1986 & n1988 ;
  assign n1990 = ~n1977 & ~n1989 ;
  assign n1991 = ~n1845 & ~n1990 ;
  assign n1992 = n1845 & n1990 ;
  assign n1993 = ~n1991 & ~n1992 ;
  assign n1994 = ~n1980 & ~n1984 ;
  assign n1995 = n1993 & ~n1994 ;
  assign n1996 = ~n1991 & ~n1995 ;
  assign n1997 = ~n1993 & n1994 ;
  assign n1998 = ~n1995 & ~n1997 ;
  assign n1999 = ~n1986 & ~n1988 ;
  assign n2000 = ~n1989 & ~n1999 ;
  assign n2001 = ~n1972 & ~n1974 ;
  assign n2002 = ~n1975 & ~n2001 ;
  assign n2003 = ~n1942 & ~n1944 ;
  assign n2004 = ~n1945 & ~n2003 ;
  assign n2005 = ~x96 & ~x256 ;
  assign n2006 = x96 & x256 ;
  assign n2007 = ~n2005 & ~n2006 ;
  assign n2008 = ~n2004 & n2007 ;
  assign n2009 = ~n2002 & n2008 ;
  assign n2010 = ~n2000 & n2009 ;
  assign n2011 = ~n1998 & n2010 ;
  assign n2012 = n1996 & n2011 ;
  assign n2013 = ~n1729 & n2012 ;
  assign n2014 = n1728 & ~n2013 ;
  assign n2015 = n571 & ~n2014 ;
  assign n2016 = ~n1728 & n2013 ;
  assign n2017 = n1723 & n1726 ;
  assign n2018 = ~n2016 & ~n2017 ;
  assign n2019 = ~n2015 & n2018 ;
  assign n2020 = ~x62 & ~x286 ;
  assign n2021 = x62 & x286 ;
  assign n2022 = ~n2020 & ~n2021 ;
  assign n2023 = ~x61 & ~x285 ;
  assign n2024 = x61 & x285 ;
  assign n2025 = ~n2023 & ~n2024 ;
  assign n2026 = n2022 & n2025 ;
  assign n2027 = ~n2022 & ~n2025 ;
  assign n2028 = ~n2026 & ~n2027 ;
  assign n2029 = ~x63 & ~x287 ;
  assign n2030 = x63 & x287 ;
  assign n2031 = ~n2029 & ~n2030 ;
  assign n2032 = ~n2028 & ~n2031 ;
  assign n2033 = n2028 & n2031 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = ~x57 & ~x281 ;
  assign n2036 = x57 & x281 ;
  assign n2037 = ~n2035 & ~n2036 ;
  assign n2038 = ~n2034 & ~n2037 ;
  assign n2039 = n2034 & n2037 ;
  assign n2040 = ~n2038 & ~n2039 ;
  assign n2041 = ~x59 & ~x283 ;
  assign n2042 = x59 & x283 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~x58 & ~x282 ;
  assign n2045 = x58 & x282 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = ~n2043 & ~n2046 ;
  assign n2048 = n2043 & n2046 ;
  assign n2049 = ~n2047 & ~n2048 ;
  assign n2050 = ~x60 & ~x284 ;
  assign n2051 = x60 & x284 ;
  assign n2052 = ~n2050 & ~n2051 ;
  assign n2053 = ~n2049 & ~n2052 ;
  assign n2054 = n2049 & n2052 ;
  assign n2055 = ~n2053 & ~n2054 ;
  assign n2056 = n2040 & ~n2055 ;
  assign n2057 = ~n2038 & ~n2056 ;
  assign n2058 = ~n2026 & ~n2033 ;
  assign n2059 = ~n2057 & n2058 ;
  assign n2060 = n2057 & ~n2058 ;
  assign n2061 = ~n2059 & ~n2060 ;
  assign n2062 = ~n2048 & ~n2054 ;
  assign n2063 = n2061 & n2062 ;
  assign n2064 = ~n2059 & ~n2063 ;
  assign n2065 = ~n2061 & ~n2062 ;
  assign n2066 = ~n2063 & ~n2065 ;
  assign n2067 = ~n2040 & n2055 ;
  assign n2068 = ~n2056 & ~n2067 ;
  assign n2069 = ~x49 & ~x273 ;
  assign n2070 = x49 & x273 ;
  assign n2071 = ~n2069 & ~n2070 ;
  assign n2072 = n2068 & ~n2071 ;
  assign n2073 = ~x55 & ~x279 ;
  assign n2074 = x55 & x279 ;
  assign n2075 = ~n2073 & ~n2074 ;
  assign n2076 = ~x54 & ~x278 ;
  assign n2077 = x54 & x278 ;
  assign n2078 = ~n2076 & ~n2077 ;
  assign n2079 = ~n2075 & ~n2078 ;
  assign n2080 = n2075 & n2078 ;
  assign n2081 = ~n2079 & ~n2080 ;
  assign n2082 = ~x56 & ~x280 ;
  assign n2083 = x56 & x280 ;
  assign n2084 = ~n2082 & ~n2083 ;
  assign n2085 = ~n2081 & ~n2084 ;
  assign n2086 = n2081 & n2084 ;
  assign n2087 = ~n2085 & ~n2086 ;
  assign n2088 = ~x50 & ~x274 ;
  assign n2089 = x50 & x274 ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2091 = ~n2087 & ~n2090 ;
  assign n2092 = n2087 & n2090 ;
  assign n2093 = ~n2091 & ~n2092 ;
  assign n2094 = ~x52 & ~x276 ;
  assign n2095 = x52 & x276 ;
  assign n2096 = ~n2094 & ~n2095 ;
  assign n2097 = ~x51 & ~x275 ;
  assign n2098 = x51 & x275 ;
  assign n2099 = ~n2097 & ~n2098 ;
  assign n2100 = ~n2096 & ~n2099 ;
  assign n2101 = n2096 & n2099 ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = ~x53 & ~x277 ;
  assign n2104 = x53 & x277 ;
  assign n2105 = ~n2103 & ~n2104 ;
  assign n2106 = ~n2102 & ~n2105 ;
  assign n2107 = n2102 & n2105 ;
  assign n2108 = ~n2106 & ~n2107 ;
  assign n2109 = n2093 & ~n2108 ;
  assign n2110 = ~n2093 & n2108 ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = ~n2068 & n2071 ;
  assign n2113 = ~n2072 & ~n2112 ;
  assign n2114 = n2111 & n2113 ;
  assign n2115 = ~n2072 & ~n2114 ;
  assign n2116 = n2066 & ~n2115 ;
  assign n2117 = ~n2091 & ~n2109 ;
  assign n2118 = ~n2080 & ~n2086 ;
  assign n2119 = ~n2117 & n2118 ;
  assign n2120 = n2117 & ~n2118 ;
  assign n2121 = ~n2119 & ~n2120 ;
  assign n2122 = ~n2101 & ~n2107 ;
  assign n2123 = n2121 & n2122 ;
  assign n2124 = ~n2121 & ~n2122 ;
  assign n2125 = ~n2123 & ~n2124 ;
  assign n2126 = ~n2066 & n2115 ;
  assign n2127 = ~n2116 & ~n2126 ;
  assign n2128 = n2125 & n2127 ;
  assign n2129 = ~n2116 & ~n2128 ;
  assign n2130 = ~n2064 & ~n2129 ;
  assign n2131 = n2064 & n2129 ;
  assign n2132 = ~n2130 & ~n2131 ;
  assign n2133 = ~n2119 & ~n2123 ;
  assign n2134 = n2132 & ~n2133 ;
  assign n2135 = ~n2130 & ~n2134 ;
  assign n2136 = ~n2132 & n2133 ;
  assign n2137 = ~n2134 & ~n2136 ;
  assign n2138 = ~n2125 & ~n2127 ;
  assign n2139 = ~n2128 & ~n2138 ;
  assign n2140 = ~n2111 & ~n2113 ;
  assign n2141 = ~n2114 & ~n2140 ;
  assign n2142 = ~x33 & ~x257 ;
  assign n2143 = x33 & x257 ;
  assign n2144 = ~n2142 & ~n2143 ;
  assign n2145 = n2141 & ~n2144 ;
  assign n2146 = ~x40 & ~x264 ;
  assign n2147 = x40 & x264 ;
  assign n2148 = ~n2146 & ~n2147 ;
  assign n2149 = ~x39 & ~x263 ;
  assign n2150 = x39 & x263 ;
  assign n2151 = ~n2149 & ~n2150 ;
  assign n2152 = ~n2148 & ~n2151 ;
  assign n2153 = n2148 & n2151 ;
  assign n2154 = ~n2152 & ~n2153 ;
  assign n2155 = ~x41 & ~x265 ;
  assign n2156 = x41 & x265 ;
  assign n2157 = ~n2155 & ~n2156 ;
  assign n2158 = ~n2154 & ~n2157 ;
  assign n2159 = n2154 & n2157 ;
  assign n2160 = ~n2158 & ~n2159 ;
  assign n2161 = ~x35 & ~x259 ;
  assign n2162 = x35 & x259 ;
  assign n2163 = ~n2161 & ~n2162 ;
  assign n2164 = ~n2160 & ~n2163 ;
  assign n2165 = n2160 & n2163 ;
  assign n2166 = ~n2164 & ~n2165 ;
  assign n2167 = ~x37 & ~x261 ;
  assign n2168 = x37 & x261 ;
  assign n2169 = ~n2167 & ~n2168 ;
  assign n2170 = ~x36 & ~x260 ;
  assign n2171 = x36 & x260 ;
  assign n2172 = ~n2170 & ~n2171 ;
  assign n2173 = ~n2169 & ~n2172 ;
  assign n2174 = n2169 & n2172 ;
  assign n2175 = ~n2173 & ~n2174 ;
  assign n2176 = ~x38 & ~x262 ;
  assign n2177 = x38 & x262 ;
  assign n2178 = ~n2176 & ~n2177 ;
  assign n2179 = ~n2175 & ~n2178 ;
  assign n2180 = n2175 & n2178 ;
  assign n2181 = ~n2179 & ~n2180 ;
  assign n2182 = n2166 & ~n2181 ;
  assign n2183 = ~n2166 & n2181 ;
  assign n2184 = ~n2182 & ~n2183 ;
  assign n2185 = ~x47 & ~x271 ;
  assign n2186 = x47 & x271 ;
  assign n2187 = ~n2185 & ~n2186 ;
  assign n2188 = ~x46 & ~x270 ;
  assign n2189 = x46 & x270 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2191 = ~n2187 & ~n2190 ;
  assign n2192 = n2187 & n2190 ;
  assign n2193 = ~n2191 & ~n2192 ;
  assign n2194 = ~x48 & ~x272 ;
  assign n2195 = x48 & x272 ;
  assign n2196 = ~n2194 & ~n2195 ;
  assign n2197 = ~n2193 & ~n2196 ;
  assign n2198 = n2193 & n2196 ;
  assign n2199 = ~n2197 & ~n2198 ;
  assign n2200 = ~x42 & ~x266 ;
  assign n2201 = x42 & x266 ;
  assign n2202 = ~n2200 & ~n2201 ;
  assign n2203 = ~n2199 & ~n2202 ;
  assign n2204 = n2199 & n2202 ;
  assign n2205 = ~n2203 & ~n2204 ;
  assign n2206 = ~x44 & ~x268 ;
  assign n2207 = x44 & x268 ;
  assign n2208 = ~n2206 & ~n2207 ;
  assign n2209 = ~x43 & ~x267 ;
  assign n2210 = x43 & x267 ;
  assign n2211 = ~n2209 & ~n2210 ;
  assign n2212 = ~n2208 & ~n2211 ;
  assign n2213 = n2208 & n2211 ;
  assign n2214 = ~n2212 & ~n2213 ;
  assign n2215 = ~x45 & ~x269 ;
  assign n2216 = x45 & x269 ;
  assign n2217 = ~n2215 & ~n2216 ;
  assign n2218 = ~n2214 & ~n2217 ;
  assign n2219 = n2214 & n2217 ;
  assign n2220 = ~n2218 & ~n2219 ;
  assign n2221 = n2205 & ~n2220 ;
  assign n2222 = ~n2205 & n2220 ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = ~x34 & ~x258 ;
  assign n2225 = x34 & x258 ;
  assign n2226 = ~n2224 & ~n2225 ;
  assign n2227 = n2223 & ~n2226 ;
  assign n2228 = ~n2223 & n2226 ;
  assign n2229 = ~n2227 & ~n2228 ;
  assign n2230 = n2184 & n2229 ;
  assign n2231 = ~n2184 & ~n2229 ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = ~n2141 & n2144 ;
  assign n2234 = ~n2145 & ~n2233 ;
  assign n2235 = n2232 & n2234 ;
  assign n2236 = ~n2145 & ~n2235 ;
  assign n2237 = n2139 & ~n2236 ;
  assign n2238 = ~n2164 & ~n2182 ;
  assign n2239 = ~n2153 & ~n2159 ;
  assign n2240 = ~n2238 & n2239 ;
  assign n2241 = n2238 & ~n2239 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2243 = ~n2174 & ~n2180 ;
  assign n2244 = n2242 & n2243 ;
  assign n2245 = ~n2242 & ~n2243 ;
  assign n2246 = ~n2244 & ~n2245 ;
  assign n2247 = ~n2203 & ~n2221 ;
  assign n2248 = ~n2192 & ~n2198 ;
  assign n2249 = ~n2247 & n2248 ;
  assign n2250 = n2247 & ~n2248 ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = ~n2213 & ~n2219 ;
  assign n2253 = n2251 & n2252 ;
  assign n2254 = ~n2251 & ~n2252 ;
  assign n2255 = ~n2253 & ~n2254 ;
  assign n2256 = ~n2227 & ~n2230 ;
  assign n2257 = n2255 & ~n2256 ;
  assign n2258 = ~n2255 & n2256 ;
  assign n2259 = ~n2257 & ~n2258 ;
  assign n2260 = n2246 & n2259 ;
  assign n2261 = ~n2246 & ~n2259 ;
  assign n2262 = ~n2260 & ~n2261 ;
  assign n2263 = ~n2139 & n2236 ;
  assign n2264 = ~n2237 & ~n2263 ;
  assign n2265 = n2262 & n2264 ;
  assign n2266 = ~n2237 & ~n2265 ;
  assign n2267 = n2137 & ~n2266 ;
  assign n2268 = ~n2249 & ~n2253 ;
  assign n2269 = ~n2257 & ~n2260 ;
  assign n2270 = ~n2268 & ~n2269 ;
  assign n2271 = n2268 & n2269 ;
  assign n2272 = ~n2270 & ~n2271 ;
  assign n2273 = ~n2240 & ~n2244 ;
  assign n2274 = n2272 & ~n2273 ;
  assign n2275 = ~n2272 & n2273 ;
  assign n2276 = ~n2274 & ~n2275 ;
  assign n2277 = ~n2137 & n2266 ;
  assign n2278 = ~n2267 & ~n2277 ;
  assign n2279 = n2276 & n2278 ;
  assign n2280 = ~n2267 & ~n2279 ;
  assign n2281 = ~n2135 & ~n2280 ;
  assign n2282 = n2135 & n2280 ;
  assign n2283 = ~n2281 & ~n2282 ;
  assign n2284 = ~n2270 & ~n2274 ;
  assign n2285 = n2283 & ~n2284 ;
  assign n2286 = ~n2281 & ~n2285 ;
  assign n2287 = ~n2283 & n2284 ;
  assign n2288 = ~n2285 & ~n2287 ;
  assign n2289 = ~n2276 & ~n2278 ;
  assign n2290 = ~n2279 & ~n2289 ;
  assign n2291 = ~n2262 & ~n2264 ;
  assign n2292 = ~n2265 & ~n2291 ;
  assign n2293 = ~n2232 & ~n2234 ;
  assign n2294 = ~n2235 & ~n2293 ;
  assign n2295 = ~x32 & ~x256 ;
  assign n2296 = x32 & x256 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2298 = ~n2294 & n2297 ;
  assign n2299 = ~n2292 & n2298 ;
  assign n2300 = ~n2290 & n2299 ;
  assign n2301 = ~n2288 & n2300 ;
  assign n2302 = n2286 & n2301 ;
  assign n2303 = ~n2019 & n2302 ;
  assign n2304 = n2016 & n2017 ;
  assign n2305 = n571 & n2304 ;
  assign n2306 = ~n2303 & n2305 ;
  assign n2307 = ~n571 & n2304 ;
  assign n2308 = n2015 & ~n2018 ;
  assign n2309 = ~n2307 & ~n2308 ;
  assign n2310 = n2303 & ~n2309 ;
  assign n2311 = ~n2306 & ~n2310 ;
  assign n2312 = ~n2303 & n2309 ;
  assign n2313 = ~x30 & ~x286 ;
  assign n2314 = x30 & x286 ;
  assign n2315 = ~n2313 & ~n2314 ;
  assign n2316 = ~x29 & ~x285 ;
  assign n2317 = x29 & x285 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = n2315 & n2318 ;
  assign n2320 = ~n2315 & ~n2318 ;
  assign n2321 = ~n2319 & ~n2320 ;
  assign n2322 = ~x31 & ~x287 ;
  assign n2323 = x31 & x287 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = ~n2321 & ~n2324 ;
  assign n2326 = n2321 & n2324 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = ~x25 & ~x281 ;
  assign n2329 = x25 & x281 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = ~n2327 & ~n2330 ;
  assign n2332 = n2327 & n2330 ;
  assign n2333 = ~n2331 & ~n2332 ;
  assign n2334 = ~x27 & ~x283 ;
  assign n2335 = x27 & x283 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = ~x26 & ~x282 ;
  assign n2338 = x26 & x282 ;
  assign n2339 = ~n2337 & ~n2338 ;
  assign n2340 = ~n2336 & ~n2339 ;
  assign n2341 = n2336 & n2339 ;
  assign n2342 = ~n2340 & ~n2341 ;
  assign n2343 = ~x28 & ~x284 ;
  assign n2344 = x28 & x284 ;
  assign n2345 = ~n2343 & ~n2344 ;
  assign n2346 = ~n2342 & ~n2345 ;
  assign n2347 = n2342 & n2345 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = n2333 & ~n2348 ;
  assign n2350 = ~n2331 & ~n2349 ;
  assign n2351 = ~n2319 & ~n2326 ;
  assign n2352 = ~n2350 & n2351 ;
  assign n2353 = n2350 & ~n2351 ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = ~n2341 & ~n2347 ;
  assign n2356 = n2354 & n2355 ;
  assign n2357 = ~n2352 & ~n2356 ;
  assign n2358 = ~n2354 & ~n2355 ;
  assign n2359 = ~n2356 & ~n2358 ;
  assign n2360 = ~n2333 & n2348 ;
  assign n2361 = ~n2349 & ~n2360 ;
  assign n2362 = ~x17 & ~x273 ;
  assign n2363 = x17 & x273 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = n2361 & ~n2364 ;
  assign n2366 = ~x23 & ~x279 ;
  assign n2367 = x23 & x279 ;
  assign n2368 = ~n2366 & ~n2367 ;
  assign n2369 = ~x22 & ~x278 ;
  assign n2370 = x22 & x278 ;
  assign n2371 = ~n2369 & ~n2370 ;
  assign n2372 = ~n2368 & ~n2371 ;
  assign n2373 = n2368 & n2371 ;
  assign n2374 = ~n2372 & ~n2373 ;
  assign n2375 = ~x24 & ~x280 ;
  assign n2376 = x24 & x280 ;
  assign n2377 = ~n2375 & ~n2376 ;
  assign n2378 = ~n2374 & ~n2377 ;
  assign n2379 = n2374 & n2377 ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = ~x18 & ~x274 ;
  assign n2382 = x18 & x274 ;
  assign n2383 = ~n2381 & ~n2382 ;
  assign n2384 = ~n2380 & ~n2383 ;
  assign n2385 = n2380 & n2383 ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2387 = ~x20 & ~x276 ;
  assign n2388 = x20 & x276 ;
  assign n2389 = ~n2387 & ~n2388 ;
  assign n2390 = ~x19 & ~x275 ;
  assign n2391 = x19 & x275 ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = ~n2389 & ~n2392 ;
  assign n2394 = n2389 & n2392 ;
  assign n2395 = ~n2393 & ~n2394 ;
  assign n2396 = ~x21 & ~x277 ;
  assign n2397 = x21 & x277 ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = ~n2395 & ~n2398 ;
  assign n2400 = n2395 & n2398 ;
  assign n2401 = ~n2399 & ~n2400 ;
  assign n2402 = n2386 & ~n2401 ;
  assign n2403 = ~n2386 & n2401 ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = ~n2361 & n2364 ;
  assign n2406 = ~n2365 & ~n2405 ;
  assign n2407 = n2404 & n2406 ;
  assign n2408 = ~n2365 & ~n2407 ;
  assign n2409 = n2359 & ~n2408 ;
  assign n2410 = ~n2384 & ~n2402 ;
  assign n2411 = ~n2373 & ~n2379 ;
  assign n2412 = ~n2410 & n2411 ;
  assign n2413 = n2410 & ~n2411 ;
  assign n2414 = ~n2412 & ~n2413 ;
  assign n2415 = ~n2394 & ~n2400 ;
  assign n2416 = n2414 & n2415 ;
  assign n2417 = ~n2414 & ~n2415 ;
  assign n2418 = ~n2416 & ~n2417 ;
  assign n2419 = ~n2359 & n2408 ;
  assign n2420 = ~n2409 & ~n2419 ;
  assign n2421 = n2418 & n2420 ;
  assign n2422 = ~n2409 & ~n2421 ;
  assign n2423 = ~n2357 & ~n2422 ;
  assign n2424 = n2357 & n2422 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = ~n2412 & ~n2416 ;
  assign n2427 = n2425 & ~n2426 ;
  assign n2428 = ~n2423 & ~n2427 ;
  assign n2429 = ~n2425 & n2426 ;
  assign n2430 = ~n2427 & ~n2429 ;
  assign n2431 = ~n2418 & ~n2420 ;
  assign n2432 = ~n2421 & ~n2431 ;
  assign n2433 = ~n2404 & ~n2406 ;
  assign n2434 = ~n2407 & ~n2433 ;
  assign n2435 = ~x1 & ~x257 ;
  assign n2436 = x1 & x257 ;
  assign n2437 = ~n2435 & ~n2436 ;
  assign n2438 = n2434 & ~n2437 ;
  assign n2439 = ~x8 & ~x264 ;
  assign n2440 = x8 & x264 ;
  assign n2441 = ~n2439 & ~n2440 ;
  assign n2442 = ~x7 & ~x263 ;
  assign n2443 = x7 & x263 ;
  assign n2444 = ~n2442 & ~n2443 ;
  assign n2445 = ~n2441 & ~n2444 ;
  assign n2446 = n2441 & n2444 ;
  assign n2447 = ~n2445 & ~n2446 ;
  assign n2448 = ~x9 & ~x265 ;
  assign n2449 = x9 & x265 ;
  assign n2450 = ~n2448 & ~n2449 ;
  assign n2451 = ~n2447 & ~n2450 ;
  assign n2452 = n2447 & n2450 ;
  assign n2453 = ~n2451 & ~n2452 ;
  assign n2454 = ~x3 & ~x259 ;
  assign n2455 = x3 & x259 ;
  assign n2456 = ~n2454 & ~n2455 ;
  assign n2457 = ~n2453 & ~n2456 ;
  assign n2458 = n2453 & n2456 ;
  assign n2459 = ~n2457 & ~n2458 ;
  assign n2460 = ~x5 & ~x261 ;
  assign n2461 = x5 & x261 ;
  assign n2462 = ~n2460 & ~n2461 ;
  assign n2463 = ~x4 & ~x260 ;
  assign n2464 = x4 & x260 ;
  assign n2465 = ~n2463 & ~n2464 ;
  assign n2466 = ~n2462 & ~n2465 ;
  assign n2467 = n2462 & n2465 ;
  assign n2468 = ~n2466 & ~n2467 ;
  assign n2469 = ~x6 & ~x262 ;
  assign n2470 = x6 & x262 ;
  assign n2471 = ~n2469 & ~n2470 ;
  assign n2472 = ~n2468 & ~n2471 ;
  assign n2473 = n2468 & n2471 ;
  assign n2474 = ~n2472 & ~n2473 ;
  assign n2475 = n2459 & ~n2474 ;
  assign n2476 = ~n2459 & n2474 ;
  assign n2477 = ~n2475 & ~n2476 ;
  assign n2478 = ~x15 & ~x271 ;
  assign n2479 = x15 & x271 ;
  assign n2480 = ~n2478 & ~n2479 ;
  assign n2481 = ~x14 & ~x270 ;
  assign n2482 = x14 & x270 ;
  assign n2483 = ~n2481 & ~n2482 ;
  assign n2484 = ~n2480 & ~n2483 ;
  assign n2485 = n2480 & n2483 ;
  assign n2486 = ~n2484 & ~n2485 ;
  assign n2487 = ~x16 & ~x272 ;
  assign n2488 = x16 & x272 ;
  assign n2489 = ~n2487 & ~n2488 ;
  assign n2490 = ~n2486 & ~n2489 ;
  assign n2491 = n2486 & n2489 ;
  assign n2492 = ~n2490 & ~n2491 ;
  assign n2493 = ~x10 & ~x266 ;
  assign n2494 = x10 & x266 ;
  assign n2495 = ~n2493 & ~n2494 ;
  assign n2496 = ~n2492 & ~n2495 ;
  assign n2497 = n2492 & n2495 ;
  assign n2498 = ~n2496 & ~n2497 ;
  assign n2499 = ~x12 & ~x268 ;
  assign n2500 = x12 & x268 ;
  assign n2501 = ~n2499 & ~n2500 ;
  assign n2502 = ~x11 & ~x267 ;
  assign n2503 = x11 & x267 ;
  assign n2504 = ~n2502 & ~n2503 ;
  assign n2505 = ~n2501 & ~n2504 ;
  assign n2506 = n2501 & n2504 ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = ~x13 & ~x269 ;
  assign n2509 = x13 & x269 ;
  assign n2510 = ~n2508 & ~n2509 ;
  assign n2511 = ~n2507 & ~n2510 ;
  assign n2512 = n2507 & n2510 ;
  assign n2513 = ~n2511 & ~n2512 ;
  assign n2514 = n2498 & ~n2513 ;
  assign n2515 = ~n2498 & n2513 ;
  assign n2516 = ~n2514 & ~n2515 ;
  assign n2517 = ~x2 & ~x258 ;
  assign n2518 = x2 & x258 ;
  assign n2519 = ~n2517 & ~n2518 ;
  assign n2520 = n2516 & ~n2519 ;
  assign n2521 = ~n2516 & n2519 ;
  assign n2522 = ~n2520 & ~n2521 ;
  assign n2523 = n2477 & n2522 ;
  assign n2524 = ~n2477 & ~n2522 ;
  assign n2525 = ~n2523 & ~n2524 ;
  assign n2526 = ~n2434 & n2437 ;
  assign n2527 = ~n2438 & ~n2526 ;
  assign n2528 = n2525 & n2527 ;
  assign n2529 = ~n2438 & ~n2528 ;
  assign n2530 = n2432 & ~n2529 ;
  assign n2531 = ~n2457 & ~n2475 ;
  assign n2532 = ~n2446 & ~n2452 ;
  assign n2533 = ~n2531 & n2532 ;
  assign n2534 = n2531 & ~n2532 ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2536 = ~n2467 & ~n2473 ;
  assign n2537 = n2535 & n2536 ;
  assign n2538 = ~n2535 & ~n2536 ;
  assign n2539 = ~n2537 & ~n2538 ;
  assign n2540 = ~n2496 & ~n2514 ;
  assign n2541 = ~n2485 & ~n2491 ;
  assign n2542 = ~n2540 & n2541 ;
  assign n2543 = n2540 & ~n2541 ;
  assign n2544 = ~n2542 & ~n2543 ;
  assign n2545 = ~n2506 & ~n2512 ;
  assign n2546 = n2544 & n2545 ;
  assign n2547 = ~n2544 & ~n2545 ;
  assign n2548 = ~n2546 & ~n2547 ;
  assign n2549 = ~n2520 & ~n2523 ;
  assign n2550 = n2548 & ~n2549 ;
  assign n2551 = ~n2548 & n2549 ;
  assign n2552 = ~n2550 & ~n2551 ;
  assign n2553 = n2539 & n2552 ;
  assign n2554 = ~n2539 & ~n2552 ;
  assign n2555 = ~n2553 & ~n2554 ;
  assign n2556 = ~n2432 & n2529 ;
  assign n2557 = ~n2530 & ~n2556 ;
  assign n2558 = n2555 & n2557 ;
  assign n2559 = ~n2530 & ~n2558 ;
  assign n2560 = n2430 & ~n2559 ;
  assign n2561 = ~n2542 & ~n2546 ;
  assign n2562 = ~n2550 & ~n2553 ;
  assign n2563 = ~n2561 & ~n2562 ;
  assign n2564 = n2561 & n2562 ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = ~n2533 & ~n2537 ;
  assign n2567 = n2565 & ~n2566 ;
  assign n2568 = ~n2565 & n2566 ;
  assign n2569 = ~n2567 & ~n2568 ;
  assign n2570 = ~n2430 & n2559 ;
  assign n2571 = ~n2560 & ~n2570 ;
  assign n2572 = n2569 & n2571 ;
  assign n2573 = ~n2560 & ~n2572 ;
  assign n2574 = ~n2428 & ~n2573 ;
  assign n2575 = n2428 & n2573 ;
  assign n2576 = ~n2574 & ~n2575 ;
  assign n2577 = ~n2563 & ~n2567 ;
  assign n2578 = n2576 & ~n2577 ;
  assign n2579 = ~n2574 & ~n2578 ;
  assign n2580 = ~n2576 & n2577 ;
  assign n2581 = ~n2578 & ~n2580 ;
  assign n2582 = ~n2555 & ~n2557 ;
  assign n2583 = ~n2558 & ~n2582 ;
  assign n2584 = ~n2525 & ~n2527 ;
  assign n2585 = ~n2528 & ~n2584 ;
  assign n2586 = ~x0 & ~x256 ;
  assign n2587 = x0 & x256 ;
  assign n2588 = ~n2586 & ~n2587 ;
  assign n2589 = ~n2585 & n2588 ;
  assign n2590 = ~n2583 & n2589 ;
  assign n2591 = ~n2569 & ~n2571 ;
  assign n2592 = ~n2572 & ~n2591 ;
  assign n2593 = n2590 & ~n2592 ;
  assign n2594 = ~n2581 & n2593 ;
  assign n2595 = n2579 & n2594 ;
  assign n2596 = ~n2312 & n2595 ;
  assign n2597 = ~n2311 & n2596 ;
  assign n2598 = n2303 & n2305 ;
  assign n2599 = ~n2597 & n2598 ;
  assign n2600 = ~n1139 & ~n1143 ;
  assign n2601 = ~n1144 & ~n2600 ;
  assign n2602 = n861 & ~n1151 ;
  assign n2603 = n1131 & ~n1149 ;
  assign n2604 = ~n1150 & ~n2603 ;
  assign n2605 = n841 & ~n859 ;
  assign n2606 = ~n860 & ~n2605 ;
  assign n2607 = n2604 & ~n2606 ;
  assign n2608 = ~n854 & ~n858 ;
  assign n2609 = ~n859 & ~n2608 ;
  assign n2610 = ~n1144 & ~n1148 ;
  assign n2611 = ~n1149 & ~n2610 ;
  assign n2612 = ~n2609 & n2611 ;
  assign n2613 = n2609 & ~n2611 ;
  assign n2614 = ~n849 & ~n853 ;
  assign n2615 = ~n854 & ~n2614 ;
  assign n2616 = n2601 & ~n2615 ;
  assign n2617 = ~n1143 & n2615 ;
  assign n2618 = ~n844 & n848 ;
  assign n2619 = ~n849 & ~n2618 ;
  assign n2620 = ~n1134 & n1138 ;
  assign n2621 = ~n1139 & ~n2620 ;
  assign n2622 = ~n2619 & n2621 ;
  assign n2623 = ~n2617 & n2622 ;
  assign n2624 = ~n2616 & ~n2623 ;
  assign n2625 = ~n2613 & ~n2624 ;
  assign n2626 = ~n2612 & ~n2625 ;
  assign n2627 = ~n2607 & n2626 ;
  assign n2628 = ~n839 & ~n860 ;
  assign n2629 = ~n861 & ~n2628 ;
  assign n2630 = ~n1129 & ~n1150 ;
  assign n2631 = ~n1151 & ~n2630 ;
  assign n2632 = n2629 & ~n2631 ;
  assign n2633 = ~n2604 & n2606 ;
  assign n2634 = ~n2632 & ~n2633 ;
  assign n2635 = ~n2627 & n2634 ;
  assign n2636 = ~n2629 & n2631 ;
  assign n2637 = ~n861 & n1151 ;
  assign n2638 = ~n2636 & ~n2637 ;
  assign n2639 = ~n2635 & n2638 ;
  assign n2640 = ~n2602 & ~n2639 ;
  assign n2641 = n2601 & ~n2640 ;
  assign n2642 = n2615 & n2640 ;
  assign n2643 = ~n2641 & ~n2642 ;
  assign n2644 = n1425 & ~n1431 ;
  assign n2645 = ~n1432 & ~n2644 ;
  assign n2646 = ~n1152 & ~n1435 ;
  assign n2647 = ~n2615 & ~n2640 ;
  assign n2648 = ~n2601 & n2640 ;
  assign n2649 = ~n2647 & ~n2648 ;
  assign n2650 = n2645 & ~n2649 ;
  assign n2651 = n1427 & ~n1430 ;
  assign n2652 = ~n1431 & ~n2651 ;
  assign n2653 = ~n2619 & ~n2640 ;
  assign n2654 = ~n2621 & n2640 ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = n2652 & ~n2655 ;
  assign n2657 = ~n2650 & ~n2656 ;
  assign n2658 = ~n2645 & n2649 ;
  assign n2659 = n1423 & ~n1432 ;
  assign n2660 = ~n1433 & ~n2659 ;
  assign n2661 = ~n2609 & ~n2640 ;
  assign n2662 = ~n2611 & n2640 ;
  assign n2663 = ~n2661 & ~n2662 ;
  assign n2664 = ~n2660 & n2663 ;
  assign n2665 = ~n2658 & ~n2664 ;
  assign n2666 = ~n2657 & n2665 ;
  assign n2667 = n2607 & ~n2640 ;
  assign n2668 = ~n2607 & ~n2633 ;
  assign n2669 = ~n2640 & ~n2668 ;
  assign n2670 = ~n2604 & ~n2669 ;
  assign n2671 = ~n2667 & ~n2670 ;
  assign n2672 = n1421 & ~n1433 ;
  assign n2673 = ~n1434 & ~n2672 ;
  assign n2674 = ~n2671 & n2673 ;
  assign n2675 = n2660 & ~n2663 ;
  assign n2676 = ~n2674 & ~n2675 ;
  assign n2677 = ~n2666 & n2676 ;
  assign n2678 = n2602 & ~n2630 ;
  assign n2679 = ~n2632 & ~n2636 ;
  assign n2680 = ~n2640 & ~n2679 ;
  assign n2681 = ~n2631 & ~n2680 ;
  assign n2682 = ~n2678 & ~n2681 ;
  assign n2683 = ~n1419 & ~n1434 ;
  assign n2684 = ~n1435 & ~n2683 ;
  assign n2685 = n2682 & ~n2684 ;
  assign n2686 = n2671 & ~n2673 ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = ~n2677 & n2687 ;
  assign n2689 = ~n2682 & n2684 ;
  assign n2690 = n1152 & n1435 ;
  assign n2691 = ~n2689 & ~n2690 ;
  assign n2692 = ~n2688 & n2691 ;
  assign n2693 = ~n2646 & ~n2692 ;
  assign n2694 = n2645 & ~n2693 ;
  assign n2695 = n2649 & n2693 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2697 = n2643 & ~n2696 ;
  assign n2698 = n2621 & ~n2640 ;
  assign n2699 = n2619 & n2640 ;
  assign n2700 = ~n2698 & ~n2699 ;
  assign n2701 = n2652 & ~n2693 ;
  assign n2702 = n2655 & n2693 ;
  assign n2703 = ~n2701 & ~n2702 ;
  assign n2704 = n2700 & ~n2703 ;
  assign n2705 = ~n2697 & ~n2704 ;
  assign n2706 = ~n2643 & n2696 ;
  assign n2707 = n2611 & ~n2640 ;
  assign n2708 = n2609 & n2640 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = n2660 & ~n2693 ;
  assign n2711 = n2663 & n2693 ;
  assign n2712 = ~n2710 & ~n2711 ;
  assign n2713 = ~n2709 & n2712 ;
  assign n2714 = ~n2706 & ~n2713 ;
  assign n2715 = ~n2705 & n2714 ;
  assign n2716 = n2606 & ~n2669 ;
  assign n2717 = ~n2667 & ~n2716 ;
  assign n2718 = n2674 & ~n2693 ;
  assign n2719 = ~n2674 & ~n2686 ;
  assign n2720 = ~n2693 & ~n2719 ;
  assign n2721 = n2671 & ~n2720 ;
  assign n2722 = ~n2718 & ~n2721 ;
  assign n2723 = n2717 & ~n2722 ;
  assign n2724 = n2709 & ~n2712 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = ~n2715 & n2725 ;
  assign n2727 = n2629 & ~n2680 ;
  assign n2728 = ~n2678 & ~n2727 ;
  assign n2729 = ~n1152 & n2689 ;
  assign n2730 = ~n2685 & ~n2689 ;
  assign n2731 = ~n2693 & ~n2730 ;
  assign n2732 = n2682 & ~n2731 ;
  assign n2733 = ~n2729 & ~n2732 ;
  assign n2734 = ~n2728 & n2733 ;
  assign n2735 = ~n2717 & n2722 ;
  assign n2736 = ~n2734 & ~n2735 ;
  assign n2737 = ~n2726 & n2736 ;
  assign n2738 = n2728 & ~n2733 ;
  assign n2739 = n1436 & ~n1437 ;
  assign n2740 = ~n2738 & ~n2739 ;
  assign n2741 = ~n2737 & n2740 ;
  assign n2742 = ~n1438 & ~n2741 ;
  assign n2743 = ~n2643 & ~n2742 ;
  assign n2744 = ~n2696 & n2742 ;
  assign n2745 = ~n2743 & ~n2744 ;
  assign n2746 = ~n1439 & ~n1724 ;
  assign n2747 = n1439 & n1724 ;
  assign n2748 = ~n1707 & ~n1722 ;
  assign n2749 = ~n1723 & ~n2748 ;
  assign n2750 = ~n2673 & ~n2720 ;
  assign n2751 = ~n2718 & ~n2750 ;
  assign n2752 = n1709 & ~n1721 ;
  assign n2753 = ~n1722 & ~n2752 ;
  assign n2754 = ~n2751 & n2753 ;
  assign n2755 = n1713 & ~n1719 ;
  assign n2756 = ~n1720 & ~n2755 ;
  assign n2757 = n2649 & ~n2693 ;
  assign n2758 = n2645 & n2693 ;
  assign n2759 = ~n2757 & ~n2758 ;
  assign n2760 = ~n2756 & ~n2759 ;
  assign n2761 = n1715 & ~n1718 ;
  assign n2762 = ~n1719 & ~n2761 ;
  assign n2763 = n2655 & ~n2693 ;
  assign n2764 = n2652 & n2693 ;
  assign n2765 = ~n2763 & ~n2764 ;
  assign n2766 = n2762 & n2765 ;
  assign n2767 = ~n2760 & n2766 ;
  assign n2768 = n2756 & n2759 ;
  assign n2769 = n1711 & ~n1720 ;
  assign n2770 = ~n1721 & ~n2769 ;
  assign n2771 = n2663 & ~n2693 ;
  assign n2772 = n2660 & n2693 ;
  assign n2773 = ~n2771 & ~n2772 ;
  assign n2774 = n2770 & n2773 ;
  assign n2775 = ~n2768 & ~n2774 ;
  assign n2776 = ~n2767 & n2775 ;
  assign n2777 = ~n2770 & ~n2773 ;
  assign n2778 = ~n2776 & ~n2777 ;
  assign n2779 = ~n2754 & ~n2778 ;
  assign n2780 = n2751 & ~n2753 ;
  assign n2781 = ~n2684 & ~n2731 ;
  assign n2782 = ~n2729 & ~n2781 ;
  assign n2783 = ~n2749 & n2782 ;
  assign n2784 = ~n1440 & ~n1723 ;
  assign n2785 = ~n2783 & ~n2784 ;
  assign n2786 = ~n2780 & n2785 ;
  assign n2787 = ~n2779 & n2786 ;
  assign n2788 = ~n1723 & n2782 ;
  assign n2789 = n1440 & ~n2748 ;
  assign n2790 = ~n2788 & n2789 ;
  assign n2791 = ~n2787 & ~n2790 ;
  assign n2792 = n2749 & n2791 ;
  assign n2793 = n2782 & ~n2791 ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2795 = n1438 & n2738 ;
  assign n2796 = ~n2734 & ~n2738 ;
  assign n2797 = ~n2742 & ~n2796 ;
  assign n2798 = n2733 & ~n2797 ;
  assign n2799 = ~n2795 & ~n2798 ;
  assign n2800 = n2794 & n2799 ;
  assign n2801 = ~n2759 & ~n2791 ;
  assign n2802 = n2756 & n2791 ;
  assign n2803 = ~n2801 & ~n2802 ;
  assign n2804 = ~n2745 & n2803 ;
  assign n2805 = ~n2762 & n2791 ;
  assign n2806 = n2765 & ~n2791 ;
  assign n2807 = ~n2805 & ~n2806 ;
  assign n2808 = n2700 & ~n2742 ;
  assign n2809 = n2703 & n2742 ;
  assign n2810 = ~n2808 & ~n2809 ;
  assign n2811 = n2807 & ~n2810 ;
  assign n2812 = ~n2804 & n2811 ;
  assign n2813 = n2745 & ~n2803 ;
  assign n2814 = n2709 & ~n2742 ;
  assign n2815 = n2712 & n2742 ;
  assign n2816 = ~n2814 & ~n2815 ;
  assign n2817 = ~n2773 & ~n2791 ;
  assign n2818 = n2770 & n2791 ;
  assign n2819 = ~n2817 & ~n2818 ;
  assign n2820 = ~n2816 & ~n2819 ;
  assign n2821 = ~n2813 & ~n2820 ;
  assign n2822 = ~n2812 & n2821 ;
  assign n2823 = n2723 & ~n2742 ;
  assign n2824 = ~n2723 & ~n2735 ;
  assign n2825 = ~n2742 & ~n2824 ;
  assign n2826 = n2722 & ~n2825 ;
  assign n2827 = ~n2823 & ~n2826 ;
  assign n2828 = n2753 & n2791 ;
  assign n2829 = n2751 & ~n2791 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = n2827 & n2830 ;
  assign n2832 = n2816 & n2819 ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2834 = ~n2822 & n2833 ;
  assign n2835 = ~n2827 & ~n2830 ;
  assign n2836 = ~n2794 & ~n2799 ;
  assign n2837 = ~n2835 & ~n2836 ;
  assign n2838 = ~n2834 & n2837 ;
  assign n2839 = ~n2800 & ~n2838 ;
  assign n2840 = ~n2747 & ~n2839 ;
  assign n2841 = ~n2746 & ~n2840 ;
  assign n2842 = ~n2745 & ~n2841 ;
  assign n2843 = ~n2803 & n2841 ;
  assign n2844 = ~n2842 & ~n2843 ;
  assign n2845 = n1998 & ~n2010 ;
  assign n2846 = ~n2011 & ~n2845 ;
  assign n2847 = ~n2830 & n2841 ;
  assign n2848 = n2827 & ~n2841 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = n2846 & n2849 ;
  assign n2851 = n2002 & ~n2008 ;
  assign n2852 = ~n2009 & ~n2851 ;
  assign n2853 = ~n2844 & ~n2852 ;
  assign n2854 = n2004 & ~n2007 ;
  assign n2855 = ~n2008 & ~n2854 ;
  assign n2856 = ~n2810 & ~n2841 ;
  assign n2857 = ~n2807 & n2841 ;
  assign n2858 = ~n2856 & ~n2857 ;
  assign n2859 = n2855 & ~n2858 ;
  assign n2860 = ~n2853 & n2859 ;
  assign n2861 = n2844 & n2852 ;
  assign n2862 = n2000 & ~n2009 ;
  assign n2863 = ~n2010 & ~n2862 ;
  assign n2864 = ~n2819 & n2841 ;
  assign n2865 = n2816 & ~n2841 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = n2863 & n2866 ;
  assign n2868 = ~n2861 & ~n2867 ;
  assign n2869 = ~n2860 & n2868 ;
  assign n2870 = ~n2863 & ~n2866 ;
  assign n2871 = ~n2869 & ~n2870 ;
  assign n2872 = ~n2850 & ~n2871 ;
  assign n2873 = ~n2846 & ~n2849 ;
  assign n2874 = ~n2794 & n2841 ;
  assign n2875 = n2799 & ~n2841 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = ~n1996 & ~n2011 ;
  assign n2878 = ~n2012 & ~n2877 ;
  assign n2879 = ~n2876 & ~n2878 ;
  assign n2880 = ~n1729 & ~n2012 ;
  assign n2881 = ~n2879 & ~n2880 ;
  assign n2882 = ~n2873 & n2881 ;
  assign n2883 = ~n2872 & n2882 ;
  assign n2884 = ~n2012 & ~n2876 ;
  assign n2885 = n1729 & ~n2877 ;
  assign n2886 = ~n2884 & n2885 ;
  assign n2887 = ~n2883 & ~n2886 ;
  assign n2888 = ~n2844 & ~n2887 ;
  assign n2889 = n2852 & n2887 ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n2891 = ~n1728 & ~n2013 ;
  assign n2892 = n1728 & n2013 ;
  assign n2893 = ~n2876 & ~n2887 ;
  assign n2894 = n2878 & n2887 ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = ~n2728 & ~n2797 ;
  assign n2897 = ~n2795 & ~n2896 ;
  assign n2898 = ~n2794 & ~n2841 ;
  assign n2899 = n2799 & n2841 ;
  assign n2900 = ~n2898 & ~n2899 ;
  assign n2901 = n2897 & ~n2900 ;
  assign n2902 = n1727 & n2901 ;
  assign n2903 = ~n2643 & n2742 ;
  assign n2904 = ~n2696 & ~n2742 ;
  assign n2905 = ~n2903 & ~n2904 ;
  assign n2906 = ~n2803 & ~n2841 ;
  assign n2907 = ~n2745 & n2841 ;
  assign n2908 = ~n2906 & ~n2907 ;
  assign n2909 = n2905 & ~n2908 ;
  assign n2910 = ~n2810 & n2841 ;
  assign n2911 = ~n2807 & ~n2841 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = ~n2700 & n2742 ;
  assign n2914 = ~n2703 & ~n2742 ;
  assign n2915 = ~n2913 & ~n2914 ;
  assign n2916 = n2912 & n2915 ;
  assign n2917 = ~n2909 & ~n2916 ;
  assign n2918 = ~n2709 & n2742 ;
  assign n2919 = ~n2712 & ~n2742 ;
  assign n2920 = ~n2918 & ~n2919 ;
  assign n2921 = ~n2819 & ~n2841 ;
  assign n2922 = n2816 & n2841 ;
  assign n2923 = ~n2921 & ~n2922 ;
  assign n2924 = ~n2920 & n2923 ;
  assign n2925 = ~n2905 & n2908 ;
  assign n2926 = ~n2924 & ~n2925 ;
  assign n2927 = ~n2917 & n2926 ;
  assign n2928 = ~n2717 & ~n2825 ;
  assign n2929 = ~n2823 & ~n2928 ;
  assign n2930 = ~n2830 & ~n2841 ;
  assign n2931 = n2827 & n2841 ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2933 = n2929 & ~n2932 ;
  assign n2934 = n2920 & ~n2923 ;
  assign n2935 = ~n2933 & ~n2934 ;
  assign n2936 = ~n2927 & n2935 ;
  assign n2937 = ~n2897 & n2900 ;
  assign n2938 = ~n2929 & n2932 ;
  assign n2939 = ~n2937 & ~n2938 ;
  assign n2940 = ~n2936 & n2939 ;
  assign n2941 = n1725 & ~n1726 ;
  assign n2942 = ~n2901 & ~n2941 ;
  assign n2943 = ~n2940 & n2942 ;
  assign n2944 = ~n1727 & ~n2943 ;
  assign n2945 = ~n2901 & ~n2937 ;
  assign n2946 = ~n2944 & ~n2945 ;
  assign n2947 = n2900 & ~n2946 ;
  assign n2948 = ~n2902 & ~n2947 ;
  assign n2949 = n2895 & n2948 ;
  assign n2950 = ~n2908 & n2944 ;
  assign n2951 = ~n2905 & ~n2944 ;
  assign n2952 = ~n2950 & ~n2951 ;
  assign n2953 = n2890 & ~n2952 ;
  assign n2954 = ~n2855 & n2887 ;
  assign n2955 = ~n2858 & ~n2887 ;
  assign n2956 = ~n2954 & ~n2955 ;
  assign n2957 = ~n2915 & ~n2944 ;
  assign n2958 = n2912 & n2944 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = n2956 & n2959 ;
  assign n2961 = ~n2953 & n2960 ;
  assign n2962 = ~n2890 & n2952 ;
  assign n2963 = ~n2920 & ~n2944 ;
  assign n2964 = ~n2923 & n2944 ;
  assign n2965 = ~n2963 & ~n2964 ;
  assign n2966 = ~n2866 & ~n2887 ;
  assign n2967 = n2863 & n2887 ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = n2965 & ~n2968 ;
  assign n2970 = ~n2962 & ~n2969 ;
  assign n2971 = ~n2961 & n2970 ;
  assign n2972 = n2933 & ~n2944 ;
  assign n2973 = n2938 & ~n2944 ;
  assign n2974 = n2932 & ~n2973 ;
  assign n2975 = ~n2972 & ~n2974 ;
  assign n2976 = ~n2849 & ~n2887 ;
  assign n2977 = n2846 & n2887 ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = n2975 & n2978 ;
  assign n2980 = ~n2965 & n2968 ;
  assign n2981 = ~n2979 & ~n2980 ;
  assign n2982 = ~n2971 & n2981 ;
  assign n2983 = ~n2975 & ~n2978 ;
  assign n2984 = ~n2895 & ~n2948 ;
  assign n2985 = ~n2983 & ~n2984 ;
  assign n2986 = ~n2982 & n2985 ;
  assign n2987 = ~n2949 & ~n2986 ;
  assign n2988 = ~n2892 & ~n2987 ;
  assign n2989 = ~n2891 & ~n2988 ;
  assign n2990 = ~n2890 & n2989 ;
  assign n2991 = ~n2952 & ~n2989 ;
  assign n2992 = ~n2990 & ~n2991 ;
  assign n2993 = n561 & ~n567 ;
  assign n2994 = ~n568 & ~n2993 ;
  assign n2995 = n2992 & n2994 ;
  assign n2996 = n563 & ~n566 ;
  assign n2997 = ~n567 & ~n2996 ;
  assign n2998 = ~n2959 & ~n2989 ;
  assign n2999 = n2956 & n2989 ;
  assign n3000 = ~n2998 & ~n2999 ;
  assign n3001 = n2997 & n3000 ;
  assign n3002 = ~n2995 & ~n3001 ;
  assign n3003 = ~n2992 & ~n2994 ;
  assign n3004 = n559 & ~n568 ;
  assign n3005 = ~n569 & ~n3004 ;
  assign n3006 = n2965 & ~n2989 ;
  assign n3007 = n2968 & n2989 ;
  assign n3008 = ~n3006 & ~n3007 ;
  assign n3009 = ~n3005 & n3008 ;
  assign n3010 = ~n3003 & ~n3009 ;
  assign n3011 = ~n3002 & n3010 ;
  assign n3012 = n3005 & ~n3008 ;
  assign n3013 = n557 & ~n569 ;
  assign n3014 = ~n570 & ~n3013 ;
  assign n3015 = ~n2978 & n2989 ;
  assign n3016 = n2975 & ~n2989 ;
  assign n3017 = ~n3015 & ~n3016 ;
  assign n3018 = n3014 & n3017 ;
  assign n3019 = ~n3012 & ~n3018 ;
  assign n3020 = ~n3011 & n3019 ;
  assign n3021 = ~n3014 & ~n3017 ;
  assign n3022 = ~n555 & ~n570 ;
  assign n3023 = ~n571 & ~n3022 ;
  assign n3024 = ~n2895 & n2989 ;
  assign n3025 = n2948 & ~n2989 ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = ~n3023 & ~n3026 ;
  assign n3028 = ~n571 & ~n2014 ;
  assign n3029 = ~n3027 & ~n3028 ;
  assign n3030 = ~n3021 & n3029 ;
  assign n3031 = ~n3020 & n3030 ;
  assign n3032 = ~n571 & ~n3026 ;
  assign n3033 = n2014 & ~n3022 ;
  assign n3034 = ~n3032 & n3033 ;
  assign n3035 = ~n3031 & ~n3034 ;
  assign n3036 = ~n2992 & ~n3035 ;
  assign n3037 = n2994 & n3035 ;
  assign n3038 = ~n3036 & ~n3037 ;
  assign n3039 = ~n2015 & ~n2018 ;
  assign n3040 = n2015 & n2018 ;
  assign n3041 = ~n3023 & n3035 ;
  assign n3042 = n3026 & ~n3035 ;
  assign n3043 = ~n3041 & ~n3042 ;
  assign n3044 = ~n2016 & n2017 ;
  assign n3045 = ~n2897 & ~n2946 ;
  assign n3046 = ~n2902 & ~n3045 ;
  assign n3047 = ~n2895 & ~n2989 ;
  assign n3048 = n2948 & n2989 ;
  assign n3049 = ~n3047 & ~n3048 ;
  assign n3050 = n3046 & ~n3049 ;
  assign n3051 = n3044 & n3050 ;
  assign n3052 = ~n2915 & n2944 ;
  assign n3053 = n2912 & ~n2944 ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = ~n2959 & n2989 ;
  assign n3056 = n2956 & ~n2989 ;
  assign n3057 = ~n3055 & ~n3056 ;
  assign n3058 = n3054 & ~n3057 ;
  assign n3059 = ~n2890 & ~n2989 ;
  assign n3060 = ~n2952 & n2989 ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3062 = ~n2908 & ~n2944 ;
  assign n3063 = ~n2905 & n2944 ;
  assign n3064 = ~n3062 & ~n3063 ;
  assign n3065 = ~n3061 & n3064 ;
  assign n3066 = ~n3058 & ~n3065 ;
  assign n3067 = ~n2920 & n2944 ;
  assign n3068 = ~n2923 & ~n2944 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = ~n2968 & ~n2989 ;
  assign n3071 = ~n2965 & n2989 ;
  assign n3072 = ~n3070 & ~n3071 ;
  assign n3073 = ~n3069 & n3072 ;
  assign n3074 = n3061 & ~n3064 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = ~n3066 & n3075 ;
  assign n3077 = ~n2929 & ~n2973 ;
  assign n3078 = ~n2972 & ~n3077 ;
  assign n3079 = ~n2978 & ~n2989 ;
  assign n3080 = n2975 & n2989 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3082 = n3078 & ~n3081 ;
  assign n3083 = n3069 & ~n3072 ;
  assign n3084 = ~n3082 & ~n3083 ;
  assign n3085 = ~n3076 & n3084 ;
  assign n3086 = ~n3046 & n3049 ;
  assign n3087 = ~n3078 & n3081 ;
  assign n3088 = ~n3086 & ~n3087 ;
  assign n3089 = ~n3085 & n3088 ;
  assign n3090 = n2016 & ~n2017 ;
  assign n3091 = ~n3050 & ~n3090 ;
  assign n3092 = ~n3089 & n3091 ;
  assign n3093 = ~n3044 & ~n3092 ;
  assign n3094 = ~n3050 & ~n3086 ;
  assign n3095 = ~n3093 & ~n3094 ;
  assign n3096 = n3049 & ~n3095 ;
  assign n3097 = ~n3051 & ~n3096 ;
  assign n3098 = ~n3043 & n3097 ;
  assign n3099 = ~n3061 & n3093 ;
  assign n3100 = ~n3064 & ~n3093 ;
  assign n3101 = ~n3099 & ~n3100 ;
  assign n3102 = n3038 & ~n3101 ;
  assign n3103 = ~n2997 & n3035 ;
  assign n3104 = n3000 & ~n3035 ;
  assign n3105 = ~n3103 & ~n3104 ;
  assign n3106 = ~n3057 & n3093 ;
  assign n3107 = ~n3054 & ~n3093 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = n3105 & n3108 ;
  assign n3110 = ~n3102 & n3109 ;
  assign n3111 = ~n3038 & n3101 ;
  assign n3112 = ~n3072 & n3093 ;
  assign n3113 = ~n3069 & ~n3093 ;
  assign n3114 = ~n3112 & ~n3113 ;
  assign n3115 = n3008 & ~n3035 ;
  assign n3116 = n3005 & n3035 ;
  assign n3117 = ~n3115 & ~n3116 ;
  assign n3118 = n3114 & ~n3117 ;
  assign n3119 = ~n3111 & ~n3118 ;
  assign n3120 = ~n3110 & n3119 ;
  assign n3121 = n3082 & ~n3093 ;
  assign n3122 = ~n3082 & ~n3087 ;
  assign n3123 = ~n3093 & ~n3122 ;
  assign n3124 = n3081 & ~n3123 ;
  assign n3125 = ~n3121 & ~n3124 ;
  assign n3126 = ~n3017 & ~n3035 ;
  assign n3127 = n3014 & n3035 ;
  assign n3128 = ~n3126 & ~n3127 ;
  assign n3129 = n3125 & n3128 ;
  assign n3130 = ~n3114 & n3117 ;
  assign n3131 = ~n3129 & ~n3130 ;
  assign n3132 = ~n3120 & n3131 ;
  assign n3133 = ~n3125 & ~n3128 ;
  assign n3134 = n3043 & ~n3097 ;
  assign n3135 = ~n3133 & ~n3134 ;
  assign n3136 = ~n3132 & n3135 ;
  assign n3137 = ~n3098 & ~n3136 ;
  assign n3138 = ~n3040 & ~n3137 ;
  assign n3139 = ~n3039 & ~n3138 ;
  assign n3140 = ~n3038 & n3139 ;
  assign n3141 = ~n3101 & ~n3139 ;
  assign n3142 = ~n3140 & ~n3141 ;
  assign n3143 = n2292 & ~n2298 ;
  assign n3144 = ~n2299 & ~n3143 ;
  assign n3145 = n3142 & n3144 ;
  assign n3146 = n2294 & ~n2297 ;
  assign n3147 = ~n2298 & ~n3146 ;
  assign n3148 = ~n3108 & ~n3139 ;
  assign n3149 = n3105 & n3139 ;
  assign n3150 = ~n3148 & ~n3149 ;
  assign n3151 = n3147 & n3150 ;
  assign n3152 = ~n3145 & ~n3151 ;
  assign n3153 = ~n3142 & ~n3144 ;
  assign n3154 = n2290 & ~n2299 ;
  assign n3155 = ~n2300 & ~n3154 ;
  assign n3156 = n3114 & ~n3139 ;
  assign n3157 = n3117 & n3139 ;
  assign n3158 = ~n3156 & ~n3157 ;
  assign n3159 = ~n3155 & n3158 ;
  assign n3160 = ~n3153 & ~n3159 ;
  assign n3161 = ~n3152 & n3160 ;
  assign n3162 = n3155 & ~n3158 ;
  assign n3163 = n2288 & ~n2300 ;
  assign n3164 = ~n2301 & ~n3163 ;
  assign n3165 = ~n3128 & n3139 ;
  assign n3166 = n3125 & ~n3139 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = n3164 & n3167 ;
  assign n3169 = ~n3162 & ~n3168 ;
  assign n3170 = ~n3161 & n3169 ;
  assign n3171 = ~n3164 & ~n3167 ;
  assign n3172 = ~n2286 & ~n2301 ;
  assign n3173 = ~n2302 & ~n3172 ;
  assign n3174 = n3097 & ~n3139 ;
  assign n3175 = n3043 & n3139 ;
  assign n3176 = ~n3174 & ~n3175 ;
  assign n3177 = ~n3173 & ~n3176 ;
  assign n3178 = ~n2019 & ~n2302 ;
  assign n3179 = ~n3177 & ~n3178 ;
  assign n3180 = ~n3171 & n3179 ;
  assign n3181 = ~n3170 & n3180 ;
  assign n3182 = ~n2302 & ~n3176 ;
  assign n3183 = n2019 & ~n3172 ;
  assign n3184 = ~n3182 & n3183 ;
  assign n3185 = ~n3181 & ~n3184 ;
  assign n3186 = ~n3142 & ~n3185 ;
  assign n3187 = n3144 & n3185 ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3189 = ~n2303 & ~n2309 ;
  assign n3190 = n2303 & n2309 ;
  assign n3191 = ~n3173 & n3185 ;
  assign n3192 = n3176 & ~n3185 ;
  assign n3193 = ~n3191 & ~n3192 ;
  assign n3194 = ~n3046 & ~n3095 ;
  assign n3195 = ~n3051 & ~n3194 ;
  assign n3196 = n3043 & ~n3139 ;
  assign n3197 = n3097 & n3139 ;
  assign n3198 = ~n3196 & ~n3197 ;
  assign n3199 = n3195 & ~n3198 ;
  assign n3200 = n2307 & n3199 ;
  assign n3201 = ~n3195 & n3198 ;
  assign n3202 = ~n3057 & ~n3093 ;
  assign n3203 = ~n3054 & n3093 ;
  assign n3204 = ~n3202 & ~n3203 ;
  assign n3205 = ~n3108 & n3139 ;
  assign n3206 = n3105 & ~n3139 ;
  assign n3207 = ~n3205 & ~n3206 ;
  assign n3208 = n3204 & ~n3207 ;
  assign n3209 = n3038 & ~n3139 ;
  assign n3210 = n3101 & n3139 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = ~n3061 & ~n3093 ;
  assign n3213 = ~n3064 & n3093 ;
  assign n3214 = ~n3212 & ~n3213 ;
  assign n3215 = n3211 & n3214 ;
  assign n3216 = ~n3208 & ~n3215 ;
  assign n3217 = ~n3072 & ~n3093 ;
  assign n3218 = ~n3069 & n3093 ;
  assign n3219 = ~n3217 & ~n3218 ;
  assign n3220 = ~n3117 & ~n3139 ;
  assign n3221 = ~n3114 & n3139 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = ~n3219 & n3222 ;
  assign n3224 = ~n3211 & ~n3214 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = ~n3216 & n3225 ;
  assign n3227 = ~n3078 & ~n3123 ;
  assign n3228 = ~n3121 & ~n3227 ;
  assign n3229 = ~n3128 & ~n3139 ;
  assign n3230 = n3125 & n3139 ;
  assign n3231 = ~n3229 & ~n3230 ;
  assign n3232 = n3228 & ~n3231 ;
  assign n3233 = n3219 & ~n3222 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3235 = ~n3226 & n3234 ;
  assign n3236 = ~n3228 & n3231 ;
  assign n3237 = ~n3201 & ~n3236 ;
  assign n3238 = ~n3235 & n3237 ;
  assign n3239 = ~n2304 & n2308 ;
  assign n3240 = ~n3199 & ~n3239 ;
  assign n3241 = ~n3238 & n3240 ;
  assign n3242 = ~n2307 & ~n3241 ;
  assign n3243 = n3201 & ~n3242 ;
  assign n3244 = n3198 & ~n3243 ;
  assign n3245 = ~n3200 & ~n3244 ;
  assign n3246 = ~n3193 & n3245 ;
  assign n3247 = ~n3214 & ~n3242 ;
  assign n3248 = n3211 & n3242 ;
  assign n3249 = ~n3247 & ~n3248 ;
  assign n3250 = n3188 & ~n3249 ;
  assign n3251 = ~n3147 & n3185 ;
  assign n3252 = n3150 & ~n3185 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = ~n3204 & ~n3242 ;
  assign n3255 = ~n3207 & n3242 ;
  assign n3256 = ~n3254 & ~n3255 ;
  assign n3257 = n3253 & n3256 ;
  assign n3258 = ~n3250 & n3257 ;
  assign n3259 = ~n3188 & n3249 ;
  assign n3260 = ~n3219 & ~n3242 ;
  assign n3261 = ~n3222 & n3242 ;
  assign n3262 = ~n3260 & ~n3261 ;
  assign n3263 = n3158 & ~n3185 ;
  assign n3264 = n3155 & n3185 ;
  assign n3265 = ~n3263 & ~n3264 ;
  assign n3266 = n3262 & ~n3265 ;
  assign n3267 = ~n3259 & ~n3266 ;
  assign n3268 = ~n3258 & n3267 ;
  assign n3269 = n3232 & ~n3242 ;
  assign n3270 = ~n3232 & ~n3236 ;
  assign n3271 = ~n3242 & ~n3270 ;
  assign n3272 = n3231 & ~n3271 ;
  assign n3273 = ~n3269 & ~n3272 ;
  assign n3274 = ~n3167 & ~n3185 ;
  assign n3275 = n3164 & n3185 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign n3277 = n3273 & n3276 ;
  assign n3278 = ~n3262 & n3265 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = ~n3268 & n3279 ;
  assign n3281 = ~n3273 & ~n3276 ;
  assign n3282 = n3193 & ~n3245 ;
  assign n3283 = ~n3281 & ~n3282 ;
  assign n3284 = ~n3280 & n3283 ;
  assign n3285 = ~n3246 & ~n3284 ;
  assign n3286 = ~n3190 & ~n3285 ;
  assign n3287 = ~n3189 & ~n3286 ;
  assign n3288 = ~n3188 & ~n3287 ;
  assign n3289 = ~n3249 & n3287 ;
  assign n3290 = ~n3288 & ~n3289 ;
  assign n3291 = ~n3207 & ~n3242 ;
  assign n3292 = ~n3204 & n3242 ;
  assign n3293 = ~n3291 & ~n3292 ;
  assign n3294 = ~n3256 & n3287 ;
  assign n3295 = n3253 & ~n3287 ;
  assign n3296 = ~n3294 & ~n3295 ;
  assign n3297 = n3293 & ~n3296 ;
  assign n3298 = ~n3214 & n3242 ;
  assign n3299 = n3211 & ~n3242 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = ~n3290 & n3300 ;
  assign n3302 = ~n3297 & ~n3301 ;
  assign n3303 = ~n3222 & ~n3242 ;
  assign n3304 = ~n3219 & n3242 ;
  assign n3305 = ~n3303 & ~n3304 ;
  assign n3306 = ~n3265 & ~n3287 ;
  assign n3307 = ~n3262 & n3287 ;
  assign n3308 = ~n3306 & ~n3307 ;
  assign n3309 = ~n3305 & n3308 ;
  assign n3310 = n3290 & ~n3300 ;
  assign n3311 = ~n3309 & ~n3310 ;
  assign n3312 = ~n3302 & n3311 ;
  assign n3313 = ~n3228 & ~n3271 ;
  assign n3314 = ~n3269 & ~n3313 ;
  assign n3315 = ~n3276 & ~n3287 ;
  assign n3316 = n3273 & n3287 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = n3314 & ~n3317 ;
  assign n3319 = n3305 & ~n3308 ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = ~n3312 & n3320 ;
  assign n3322 = ~n3314 & n3317 ;
  assign n3323 = ~n3195 & ~n3243 ;
  assign n3324 = ~n3200 & ~n3323 ;
  assign n3325 = n3193 & ~n3287 ;
  assign n3326 = n3245 & n3287 ;
  assign n3327 = ~n3325 & ~n3326 ;
  assign n3328 = ~n3324 & n3327 ;
  assign n3329 = ~n3322 & ~n3328 ;
  assign n3330 = ~n3321 & n3329 ;
  assign n3331 = n3324 & ~n3327 ;
  assign n3332 = ~n2305 & n2310 ;
  assign n3333 = ~n3331 & ~n3332 ;
  assign n3334 = ~n3330 & n3333 ;
  assign n3335 = ~n2306 & ~n3334 ;
  assign n3336 = n3290 & ~n3335 ;
  assign n3337 = n3300 & n3335 ;
  assign n3338 = ~n3336 & ~n3337 ;
  assign n3339 = ~n3188 & n3287 ;
  assign n3340 = ~n3249 & ~n3287 ;
  assign n3341 = ~n3339 & ~n3340 ;
  assign n3342 = n2583 & ~n2589 ;
  assign n3343 = ~n2590 & ~n3342 ;
  assign n3344 = n3341 & n3343 ;
  assign n3345 = n2585 & ~n2588 ;
  assign n3346 = ~n2589 & ~n3345 ;
  assign n3347 = ~n3256 & ~n3287 ;
  assign n3348 = n3253 & n3287 ;
  assign n3349 = ~n3347 & ~n3348 ;
  assign n3350 = n3346 & n3349 ;
  assign n3351 = ~n3344 & ~n3350 ;
  assign n3352 = ~n3341 & ~n3343 ;
  assign n3353 = ~n2590 & n2592 ;
  assign n3354 = ~n2593 & ~n3353 ;
  assign n3355 = n3262 & ~n3287 ;
  assign n3356 = n3265 & n3287 ;
  assign n3357 = ~n3355 & ~n3356 ;
  assign n3358 = ~n3354 & n3357 ;
  assign n3359 = ~n3352 & ~n3358 ;
  assign n3360 = ~n3351 & n3359 ;
  assign n3361 = n3354 & ~n3357 ;
  assign n3362 = n2581 & ~n2593 ;
  assign n3363 = ~n2594 & ~n3362 ;
  assign n3364 = ~n3276 & n3287 ;
  assign n3365 = n3273 & ~n3287 ;
  assign n3366 = ~n3364 & ~n3365 ;
  assign n3367 = n3363 & n3366 ;
  assign n3368 = ~n3361 & ~n3367 ;
  assign n3369 = ~n3360 & n3368 ;
  assign n3370 = ~n3363 & ~n3366 ;
  assign n3371 = ~n2579 & ~n2594 ;
  assign n3372 = ~n2595 & ~n3371 ;
  assign n3373 = n3245 & ~n3287 ;
  assign n3374 = n3193 & n3287 ;
  assign n3375 = ~n3373 & ~n3374 ;
  assign n3376 = ~n3372 & ~n3375 ;
  assign n3377 = ~n2312 & ~n2595 ;
  assign n3378 = ~n3376 & ~n3377 ;
  assign n3379 = ~n3370 & n3378 ;
  assign n3380 = ~n3369 & n3379 ;
  assign n3381 = ~n2595 & ~n3375 ;
  assign n3382 = n2312 & ~n3371 ;
  assign n3383 = ~n3381 & n3382 ;
  assign n3384 = ~n3380 & ~n3383 ;
  assign n3385 = ~n3341 & ~n3384 ;
  assign n3386 = n3343 & n3384 ;
  assign n3387 = ~n3385 & ~n3386 ;
  assign n3388 = ~n2311 & ~n2596 ;
  assign n3389 = n2311 & n2596 ;
  assign n3390 = n2306 & n3331 ;
  assign n3391 = ~n3328 & ~n3331 ;
  assign n3392 = ~n3335 & ~n3391 ;
  assign n3393 = n3327 & ~n3392 ;
  assign n3394 = ~n3390 & ~n3393 ;
  assign n3395 = ~n3372 & n3384 ;
  assign n3396 = n3375 & ~n3384 ;
  assign n3397 = ~n3395 & ~n3396 ;
  assign n3398 = n3394 & ~n3397 ;
  assign n3399 = ~n3290 & n3335 ;
  assign n3400 = ~n3300 & ~n3335 ;
  assign n3401 = ~n3399 & ~n3400 ;
  assign n3402 = n3387 & ~n3401 ;
  assign n3403 = ~n3346 & n3384 ;
  assign n3404 = n3349 & ~n3384 ;
  assign n3405 = ~n3403 & ~n3404 ;
  assign n3406 = ~n3293 & ~n3335 ;
  assign n3407 = ~n3296 & n3335 ;
  assign n3408 = ~n3406 & ~n3407 ;
  assign n3409 = n3405 & n3408 ;
  assign n3410 = ~n3402 & n3409 ;
  assign n3411 = ~n3305 & ~n3335 ;
  assign n3412 = ~n3308 & n3335 ;
  assign n3413 = ~n3411 & ~n3412 ;
  assign n3414 = n3357 & ~n3384 ;
  assign n3415 = n3354 & n3384 ;
  assign n3416 = ~n3414 & ~n3415 ;
  assign n3417 = n3413 & ~n3416 ;
  assign n3418 = ~n3387 & n3401 ;
  assign n3419 = ~n3417 & ~n3418 ;
  assign n3420 = ~n3410 & n3419 ;
  assign n3421 = ~n3318 & ~n3322 ;
  assign n3422 = ~n3335 & ~n3421 ;
  assign n3423 = n3317 & ~n3422 ;
  assign n3424 = n3318 & ~n3335 ;
  assign n3425 = ~n3423 & ~n3424 ;
  assign n3426 = ~n3366 & ~n3384 ;
  assign n3427 = n3363 & n3384 ;
  assign n3428 = ~n3426 & ~n3427 ;
  assign n3429 = n3425 & n3428 ;
  assign n3430 = ~n3413 & n3416 ;
  assign n3431 = ~n3429 & ~n3430 ;
  assign n3432 = ~n3420 & n3431 ;
  assign n3433 = ~n3394 & n3397 ;
  assign n3434 = ~n3425 & ~n3428 ;
  assign n3435 = ~n3433 & ~n3434 ;
  assign n3436 = ~n3432 & n3435 ;
  assign n3437 = ~n3398 & ~n3436 ;
  assign n3438 = ~n3389 & ~n3437 ;
  assign n3439 = ~n3388 & ~n3438 ;
  assign n3440 = ~n3387 & ~n3439 ;
  assign n3441 = ~n3401 & n3439 ;
  assign n3442 = ~n3440 & ~n3441 ;
  assign n3443 = ~n3338 & ~n3442 ;
  assign n3444 = n3408 & n3439 ;
  assign n3445 = ~n3405 & ~n3439 ;
  assign n3446 = n3293 & n3335 ;
  assign n3447 = n3296 & ~n3335 ;
  assign n3448 = ~n3446 & ~n3447 ;
  assign n3449 = ~n3445 & ~n3448 ;
  assign n3450 = ~n3444 & n3449 ;
  assign n3451 = ~n3443 & ~n3450 ;
  assign n3452 = n3338 & n3442 ;
  assign n3453 = ~n3305 & n3335 ;
  assign n3454 = ~n3308 & ~n3335 ;
  assign n3455 = ~n3453 & ~n3454 ;
  assign n3456 = ~n3413 & n3439 ;
  assign n3457 = ~n3416 & ~n3439 ;
  assign n3458 = ~n3456 & ~n3457 ;
  assign n3459 = ~n3455 & n3458 ;
  assign n3460 = ~n3452 & ~n3459 ;
  assign n3461 = ~n3451 & n3460 ;
  assign n3462 = n3455 & ~n3458 ;
  assign n3463 = ~n3314 & ~n3422 ;
  assign n3464 = ~n3424 & ~n3463 ;
  assign n3465 = ~n3428 & ~n3439 ;
  assign n3466 = n3425 & n3439 ;
  assign n3467 = ~n3465 & ~n3466 ;
  assign n3468 = n3464 & ~n3467 ;
  assign n3469 = ~n3462 & ~n3468 ;
  assign n3470 = ~n3461 & n3469 ;
  assign n3471 = ~n3464 & n3467 ;
  assign n3472 = ~n3470 & ~n3471 ;
  assign n3473 = n3394 & n3439 ;
  assign n3474 = n3397 & ~n3439 ;
  assign n3475 = ~n3473 & ~n3474 ;
  assign n3476 = ~n3472 & n3475 ;
  assign n3477 = ~n3324 & ~n3392 ;
  assign n3478 = ~n3390 & ~n3477 ;
  assign n3479 = ~n3476 & n3478 ;
  assign n3480 = n2597 & ~n2598 ;
  assign n3481 = n3472 & ~n3475 ;
  assign n3482 = ~n3480 & ~n3481 ;
  assign n3483 = ~n3479 & n3482 ;
  assign n3484 = ~n2599 & ~n3483 ;
  assign n3485 = x224 & ~n2640 ;
  assign n3486 = x192 & n2640 ;
  assign n3487 = ~n3485 & ~n3486 ;
  assign n3488 = n2693 & ~n3487 ;
  assign n3489 = x160 & ~n2693 ;
  assign n3490 = ~n3488 & ~n3489 ;
  assign n3491 = ~n2742 & ~n3490 ;
  assign n3492 = x192 & ~n2640 ;
  assign n3493 = x224 & n2640 ;
  assign n3494 = ~n3492 & ~n3493 ;
  assign n3495 = n2742 & ~n3494 ;
  assign n3496 = ~n3491 & ~n3495 ;
  assign n3497 = n2944 & ~n3496 ;
  assign n3498 = n2742 & ~n3490 ;
  assign n3499 = ~n2742 & ~n3494 ;
  assign n3500 = ~n3498 & ~n3499 ;
  assign n3501 = n2841 & ~n3500 ;
  assign n3502 = ~n2693 & ~n3487 ;
  assign n3503 = x160 & n2693 ;
  assign n3504 = ~n3502 & ~n3503 ;
  assign n3505 = ~n2791 & ~n3504 ;
  assign n3506 = x128 & n2791 ;
  assign n3507 = ~n3505 & ~n3506 ;
  assign n3508 = ~n2841 & ~n3507 ;
  assign n3509 = ~n3501 & ~n3508 ;
  assign n3510 = ~n2944 & ~n3509 ;
  assign n3511 = ~n3497 & ~n3510 ;
  assign n3512 = n3093 & ~n3511 ;
  assign n3513 = ~n2944 & ~n3496 ;
  assign n3514 = n2944 & ~n3509 ;
  assign n3515 = ~n3513 & ~n3514 ;
  assign n3516 = n2989 & ~n3515 ;
  assign n3517 = ~n2841 & ~n3500 ;
  assign n3518 = n2841 & ~n3507 ;
  assign n3519 = ~n3517 & ~n3518 ;
  assign n3520 = ~n2887 & ~n3519 ;
  assign n3521 = x96 & n2887 ;
  assign n3522 = ~n3520 & ~n3521 ;
  assign n3523 = ~n2989 & ~n3522 ;
  assign n3524 = ~n3516 & ~n3523 ;
  assign n3525 = ~n3093 & ~n3524 ;
  assign n3526 = ~n3512 & ~n3525 ;
  assign n3527 = ~n3242 & ~n3526 ;
  assign n3528 = ~n3093 & ~n3511 ;
  assign n3529 = n3093 & ~n3524 ;
  assign n3530 = ~n3528 & ~n3529 ;
  assign n3531 = n3139 & ~n3530 ;
  assign n3532 = n2989 & ~n3522 ;
  assign n3533 = ~n2989 & ~n3515 ;
  assign n3534 = ~n3532 & ~n3533 ;
  assign n3535 = ~n3035 & ~n3534 ;
  assign n3536 = x64 & n3035 ;
  assign n3537 = ~n3535 & ~n3536 ;
  assign n3538 = ~n3139 & ~n3537 ;
  assign n3539 = ~n3531 & ~n3538 ;
  assign n3540 = n3242 & ~n3539 ;
  assign n3541 = ~n3527 & ~n3540 ;
  assign n3542 = ~n3287 & ~n3541 ;
  assign n3543 = n3139 & ~n3537 ;
  assign n3544 = ~n3139 & ~n3530 ;
  assign n3545 = ~n3543 & ~n3544 ;
  assign n3546 = ~n3185 & ~n3545 ;
  assign n3547 = x32 & n3185 ;
  assign n3548 = ~n3546 & ~n3547 ;
  assign n3549 = n3287 & ~n3548 ;
  assign n3550 = ~n3542 & ~n3549 ;
  assign n3551 = ~n3384 & ~n3550 ;
  assign n3552 = x0 & n3384 ;
  assign n3553 = ~n3551 & ~n3552 ;
  assign n3554 = ~n3439 & ~n3553 ;
  assign n3555 = ~n3287 & ~n3548 ;
  assign n3556 = n3287 & ~n3541 ;
  assign n3557 = ~n3555 & ~n3556 ;
  assign n3558 = n3335 & ~n3557 ;
  assign n3559 = n3242 & ~n3526 ;
  assign n3560 = ~n3242 & ~n3539 ;
  assign n3561 = ~n3559 & ~n3560 ;
  assign n3562 = ~n3335 & ~n3561 ;
  assign n3563 = ~n3558 & ~n3562 ;
  assign n3564 = n3439 & ~n3563 ;
  assign n3565 = ~n3554 & ~n3564 ;
  assign n3566 = ~n3484 & ~n3565 ;
  assign n3567 = ~n3335 & ~n3557 ;
  assign n3568 = n3335 & ~n3561 ;
  assign n3569 = ~n3567 & ~n3568 ;
  assign n3570 = n3484 & ~n3569 ;
  assign n3571 = ~n3566 & ~n3570 ;
  assign n3572 = x225 & ~n2640 ;
  assign n3573 = x193 & n2640 ;
  assign n3574 = ~n3572 & ~n3573 ;
  assign n3575 = n2693 & ~n3574 ;
  assign n3576 = x161 & ~n2693 ;
  assign n3577 = ~n3575 & ~n3576 ;
  assign n3578 = n2742 & ~n3577 ;
  assign n3579 = x193 & ~n2640 ;
  assign n3580 = x225 & n2640 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = ~n2742 & ~n3581 ;
  assign n3583 = ~n3578 & ~n3582 ;
  assign n3584 = ~n2841 & ~n3583 ;
  assign n3585 = ~n2693 & ~n3574 ;
  assign n3586 = x161 & n2693 ;
  assign n3587 = ~n3585 & ~n3586 ;
  assign n3588 = ~n2791 & ~n3587 ;
  assign n3589 = x129 & n2791 ;
  assign n3590 = ~n3588 & ~n3589 ;
  assign n3591 = n2841 & ~n3590 ;
  assign n3592 = ~n3584 & ~n3591 ;
  assign n3593 = ~n2887 & ~n3592 ;
  assign n3594 = x97 & n2887 ;
  assign n3595 = ~n3593 & ~n3594 ;
  assign n3596 = n2989 & ~n3595 ;
  assign n3597 = n2841 & ~n3583 ;
  assign n3598 = ~n2841 & ~n3590 ;
  assign n3599 = ~n3597 & ~n3598 ;
  assign n3600 = n2944 & ~n3599 ;
  assign n3601 = n2742 & ~n3581 ;
  assign n3602 = ~n2742 & ~n3577 ;
  assign n3603 = ~n3601 & ~n3602 ;
  assign n3604 = ~n2944 & ~n3603 ;
  assign n3605 = ~n3600 & ~n3604 ;
  assign n3606 = ~n2989 & ~n3605 ;
  assign n3607 = ~n3596 & ~n3606 ;
  assign n3608 = ~n3035 & ~n3607 ;
  assign n3609 = x65 & n3035 ;
  assign n3610 = ~n3608 & ~n3609 ;
  assign n3611 = n3139 & ~n3610 ;
  assign n3612 = n2944 & ~n3603 ;
  assign n3613 = ~n2944 & ~n3599 ;
  assign n3614 = ~n3612 & ~n3613 ;
  assign n3615 = ~n3093 & ~n3614 ;
  assign n3616 = n2989 & ~n3605 ;
  assign n3617 = ~n2989 & ~n3595 ;
  assign n3618 = ~n3616 & ~n3617 ;
  assign n3619 = n3093 & ~n3618 ;
  assign n3620 = ~n3615 & ~n3619 ;
  assign n3621 = ~n3139 & ~n3620 ;
  assign n3622 = ~n3611 & ~n3621 ;
  assign n3623 = ~n3185 & ~n3622 ;
  assign n3624 = x33 & n3185 ;
  assign n3625 = ~n3623 & ~n3624 ;
  assign n3626 = ~n3287 & ~n3625 ;
  assign n3627 = n3093 & ~n3614 ;
  assign n3628 = ~n3093 & ~n3618 ;
  assign n3629 = ~n3627 & ~n3628 ;
  assign n3630 = ~n3242 & ~n3629 ;
  assign n3631 = n3139 & ~n3620 ;
  assign n3632 = ~n3139 & ~n3610 ;
  assign n3633 = ~n3631 & ~n3632 ;
  assign n3634 = n3242 & ~n3633 ;
  assign n3635 = ~n3630 & ~n3634 ;
  assign n3636 = n3287 & ~n3635 ;
  assign n3637 = ~n3626 & ~n3636 ;
  assign n3638 = ~n3335 & ~n3637 ;
  assign n3639 = n3242 & ~n3629 ;
  assign n3640 = ~n3242 & ~n3633 ;
  assign n3641 = ~n3639 & ~n3640 ;
  assign n3642 = n3335 & ~n3641 ;
  assign n3643 = ~n3638 & ~n3642 ;
  assign n3644 = n3484 & ~n3643 ;
  assign n3645 = n3335 & ~n3637 ;
  assign n3646 = ~n3335 & ~n3641 ;
  assign n3647 = ~n3645 & ~n3646 ;
  assign n3648 = n3439 & ~n3647 ;
  assign n3649 = ~n3287 & ~n3635 ;
  assign n3650 = n3287 & ~n3625 ;
  assign n3651 = ~n3649 & ~n3650 ;
  assign n3652 = ~n3384 & ~n3651 ;
  assign n3653 = x1 & n3384 ;
  assign n3654 = ~n3652 & ~n3653 ;
  assign n3655 = ~n3439 & ~n3654 ;
  assign n3656 = ~n3648 & ~n3655 ;
  assign n3657 = ~n3484 & ~n3656 ;
  assign n3658 = ~n3644 & ~n3657 ;
  assign n3659 = x226 & ~n2640 ;
  assign n3660 = x194 & n2640 ;
  assign n3661 = ~n3659 & ~n3660 ;
  assign n3662 = n2693 & ~n3661 ;
  assign n3663 = x162 & ~n2693 ;
  assign n3664 = ~n3662 & ~n3663 ;
  assign n3665 = n2742 & ~n3664 ;
  assign n3666 = x194 & ~n2640 ;
  assign n3667 = x226 & n2640 ;
  assign n3668 = ~n3666 & ~n3667 ;
  assign n3669 = ~n2742 & ~n3668 ;
  assign n3670 = ~n3665 & ~n3669 ;
  assign n3671 = ~n2841 & ~n3670 ;
  assign n3672 = ~n2693 & ~n3661 ;
  assign n3673 = x162 & n2693 ;
  assign n3674 = ~n3672 & ~n3673 ;
  assign n3675 = ~n2791 & ~n3674 ;
  assign n3676 = x130 & n2791 ;
  assign n3677 = ~n3675 & ~n3676 ;
  assign n3678 = n2841 & ~n3677 ;
  assign n3679 = ~n3671 & ~n3678 ;
  assign n3680 = ~n2887 & ~n3679 ;
  assign n3681 = x98 & n2887 ;
  assign n3682 = ~n3680 & ~n3681 ;
  assign n3683 = n2989 & ~n3682 ;
  assign n3684 = n2841 & ~n3670 ;
  assign n3685 = ~n2841 & ~n3677 ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = n2944 & ~n3686 ;
  assign n3688 = n2742 & ~n3668 ;
  assign n3689 = ~n2742 & ~n3664 ;
  assign n3690 = ~n3688 & ~n3689 ;
  assign n3691 = ~n2944 & ~n3690 ;
  assign n3692 = ~n3687 & ~n3691 ;
  assign n3693 = ~n2989 & ~n3692 ;
  assign n3694 = ~n3683 & ~n3693 ;
  assign n3695 = ~n3035 & ~n3694 ;
  assign n3696 = x66 & n3035 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3698 = n3139 & ~n3697 ;
  assign n3699 = n2944 & ~n3690 ;
  assign n3700 = ~n2944 & ~n3686 ;
  assign n3701 = ~n3699 & ~n3700 ;
  assign n3702 = ~n3093 & ~n3701 ;
  assign n3703 = n2989 & ~n3692 ;
  assign n3704 = ~n2989 & ~n3682 ;
  assign n3705 = ~n3703 & ~n3704 ;
  assign n3706 = n3093 & ~n3705 ;
  assign n3707 = ~n3702 & ~n3706 ;
  assign n3708 = ~n3139 & ~n3707 ;
  assign n3709 = ~n3698 & ~n3708 ;
  assign n3710 = ~n3185 & ~n3709 ;
  assign n3711 = x34 & n3185 ;
  assign n3712 = ~n3710 & ~n3711 ;
  assign n3713 = ~n3287 & ~n3712 ;
  assign n3714 = n3093 & ~n3701 ;
  assign n3715 = ~n3093 & ~n3705 ;
  assign n3716 = ~n3714 & ~n3715 ;
  assign n3717 = ~n3242 & ~n3716 ;
  assign n3718 = n3139 & ~n3707 ;
  assign n3719 = ~n3139 & ~n3697 ;
  assign n3720 = ~n3718 & ~n3719 ;
  assign n3721 = n3242 & ~n3720 ;
  assign n3722 = ~n3717 & ~n3721 ;
  assign n3723 = n3287 & ~n3722 ;
  assign n3724 = ~n3713 & ~n3723 ;
  assign n3725 = ~n3335 & ~n3724 ;
  assign n3726 = n3242 & ~n3716 ;
  assign n3727 = ~n3242 & ~n3720 ;
  assign n3728 = ~n3726 & ~n3727 ;
  assign n3729 = n3335 & ~n3728 ;
  assign n3730 = ~n3725 & ~n3729 ;
  assign n3731 = n3484 & ~n3730 ;
  assign n3732 = n3335 & ~n3724 ;
  assign n3733 = ~n3335 & ~n3728 ;
  assign n3734 = ~n3732 & ~n3733 ;
  assign n3735 = n3439 & ~n3734 ;
  assign n3736 = ~n3287 & ~n3722 ;
  assign n3737 = n3287 & ~n3712 ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = ~n3384 & ~n3738 ;
  assign n3740 = x2 & n3384 ;
  assign n3741 = ~n3739 & ~n3740 ;
  assign n3742 = ~n3439 & ~n3741 ;
  assign n3743 = ~n3735 & ~n3742 ;
  assign n3744 = ~n3484 & ~n3743 ;
  assign n3745 = ~n3731 & ~n3744 ;
  assign n3746 = x227 & ~n2640 ;
  assign n3747 = x195 & n2640 ;
  assign n3748 = ~n3746 & ~n3747 ;
  assign n3749 = n2693 & ~n3748 ;
  assign n3750 = x163 & ~n2693 ;
  assign n3751 = ~n3749 & ~n3750 ;
  assign n3752 = n2742 & ~n3751 ;
  assign n3753 = x195 & ~n2640 ;
  assign n3754 = x227 & n2640 ;
  assign n3755 = ~n3753 & ~n3754 ;
  assign n3756 = ~n2742 & ~n3755 ;
  assign n3757 = ~n3752 & ~n3756 ;
  assign n3758 = ~n2841 & ~n3757 ;
  assign n3759 = ~n2693 & ~n3748 ;
  assign n3760 = x163 & n2693 ;
  assign n3761 = ~n3759 & ~n3760 ;
  assign n3762 = ~n2791 & ~n3761 ;
  assign n3763 = x131 & n2791 ;
  assign n3764 = ~n3762 & ~n3763 ;
  assign n3765 = n2841 & ~n3764 ;
  assign n3766 = ~n3758 & ~n3765 ;
  assign n3767 = ~n2887 & ~n3766 ;
  assign n3768 = x99 & n2887 ;
  assign n3769 = ~n3767 & ~n3768 ;
  assign n3770 = n2989 & ~n3769 ;
  assign n3771 = n2841 & ~n3757 ;
  assign n3772 = ~n2841 & ~n3764 ;
  assign n3773 = ~n3771 & ~n3772 ;
  assign n3774 = n2944 & ~n3773 ;
  assign n3775 = n2742 & ~n3755 ;
  assign n3776 = ~n2742 & ~n3751 ;
  assign n3777 = ~n3775 & ~n3776 ;
  assign n3778 = ~n2944 & ~n3777 ;
  assign n3779 = ~n3774 & ~n3778 ;
  assign n3780 = ~n2989 & ~n3779 ;
  assign n3781 = ~n3770 & ~n3780 ;
  assign n3782 = ~n3035 & ~n3781 ;
  assign n3783 = x67 & n3035 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = n3139 & ~n3784 ;
  assign n3786 = n2944 & ~n3777 ;
  assign n3787 = ~n2944 & ~n3773 ;
  assign n3788 = ~n3786 & ~n3787 ;
  assign n3789 = ~n3093 & ~n3788 ;
  assign n3790 = n2989 & ~n3779 ;
  assign n3791 = ~n2989 & ~n3769 ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3793 = n3093 & ~n3792 ;
  assign n3794 = ~n3789 & ~n3793 ;
  assign n3795 = ~n3139 & ~n3794 ;
  assign n3796 = ~n3785 & ~n3795 ;
  assign n3797 = ~n3185 & ~n3796 ;
  assign n3798 = x35 & n3185 ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = ~n3287 & ~n3799 ;
  assign n3801 = n3093 & ~n3788 ;
  assign n3802 = ~n3093 & ~n3792 ;
  assign n3803 = ~n3801 & ~n3802 ;
  assign n3804 = ~n3242 & ~n3803 ;
  assign n3805 = n3139 & ~n3794 ;
  assign n3806 = ~n3139 & ~n3784 ;
  assign n3807 = ~n3805 & ~n3806 ;
  assign n3808 = n3242 & ~n3807 ;
  assign n3809 = ~n3804 & ~n3808 ;
  assign n3810 = n3287 & ~n3809 ;
  assign n3811 = ~n3800 & ~n3810 ;
  assign n3812 = ~n3335 & ~n3811 ;
  assign n3813 = n3242 & ~n3803 ;
  assign n3814 = ~n3242 & ~n3807 ;
  assign n3815 = ~n3813 & ~n3814 ;
  assign n3816 = n3335 & ~n3815 ;
  assign n3817 = ~n3812 & ~n3816 ;
  assign n3818 = n3484 & ~n3817 ;
  assign n3819 = n3335 & ~n3811 ;
  assign n3820 = ~n3335 & ~n3815 ;
  assign n3821 = ~n3819 & ~n3820 ;
  assign n3822 = n3439 & ~n3821 ;
  assign n3823 = ~n3287 & ~n3809 ;
  assign n3824 = n3287 & ~n3799 ;
  assign n3825 = ~n3823 & ~n3824 ;
  assign n3826 = ~n3384 & ~n3825 ;
  assign n3827 = x3 & n3384 ;
  assign n3828 = ~n3826 & ~n3827 ;
  assign n3829 = ~n3439 & ~n3828 ;
  assign n3830 = ~n3822 & ~n3829 ;
  assign n3831 = ~n3484 & ~n3830 ;
  assign n3832 = ~n3818 & ~n3831 ;
  assign n3833 = x228 & ~n2640 ;
  assign n3834 = x196 & n2640 ;
  assign n3835 = ~n3833 & ~n3834 ;
  assign n3836 = n2693 & ~n3835 ;
  assign n3837 = x164 & ~n2693 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = n2742 & ~n3838 ;
  assign n3840 = x196 & ~n2640 ;
  assign n3841 = x228 & n2640 ;
  assign n3842 = ~n3840 & ~n3841 ;
  assign n3843 = ~n2742 & ~n3842 ;
  assign n3844 = ~n3839 & ~n3843 ;
  assign n3845 = ~n2841 & ~n3844 ;
  assign n3846 = ~n2693 & ~n3835 ;
  assign n3847 = x164 & n2693 ;
  assign n3848 = ~n3846 & ~n3847 ;
  assign n3849 = ~n2791 & ~n3848 ;
  assign n3850 = x132 & n2791 ;
  assign n3851 = ~n3849 & ~n3850 ;
  assign n3852 = n2841 & ~n3851 ;
  assign n3853 = ~n3845 & ~n3852 ;
  assign n3854 = ~n2887 & ~n3853 ;
  assign n3855 = x100 & n2887 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = n2989 & ~n3856 ;
  assign n3858 = n2841 & ~n3844 ;
  assign n3859 = ~n2841 & ~n3851 ;
  assign n3860 = ~n3858 & ~n3859 ;
  assign n3861 = n2944 & ~n3860 ;
  assign n3862 = n2742 & ~n3842 ;
  assign n3863 = ~n2742 & ~n3838 ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = ~n2944 & ~n3864 ;
  assign n3866 = ~n3861 & ~n3865 ;
  assign n3867 = ~n2989 & ~n3866 ;
  assign n3868 = ~n3857 & ~n3867 ;
  assign n3869 = ~n3035 & ~n3868 ;
  assign n3870 = x68 & n3035 ;
  assign n3871 = ~n3869 & ~n3870 ;
  assign n3872 = n3139 & ~n3871 ;
  assign n3873 = n2944 & ~n3864 ;
  assign n3874 = ~n2944 & ~n3860 ;
  assign n3875 = ~n3873 & ~n3874 ;
  assign n3876 = ~n3093 & ~n3875 ;
  assign n3877 = n2989 & ~n3866 ;
  assign n3878 = ~n2989 & ~n3856 ;
  assign n3879 = ~n3877 & ~n3878 ;
  assign n3880 = n3093 & ~n3879 ;
  assign n3881 = ~n3876 & ~n3880 ;
  assign n3882 = ~n3139 & ~n3881 ;
  assign n3883 = ~n3872 & ~n3882 ;
  assign n3884 = ~n3185 & ~n3883 ;
  assign n3885 = x36 & n3185 ;
  assign n3886 = ~n3884 & ~n3885 ;
  assign n3887 = ~n3287 & ~n3886 ;
  assign n3888 = n3093 & ~n3875 ;
  assign n3889 = ~n3093 & ~n3879 ;
  assign n3890 = ~n3888 & ~n3889 ;
  assign n3891 = ~n3242 & ~n3890 ;
  assign n3892 = n3139 & ~n3881 ;
  assign n3893 = ~n3139 & ~n3871 ;
  assign n3894 = ~n3892 & ~n3893 ;
  assign n3895 = n3242 & ~n3894 ;
  assign n3896 = ~n3891 & ~n3895 ;
  assign n3897 = n3287 & ~n3896 ;
  assign n3898 = ~n3887 & ~n3897 ;
  assign n3899 = ~n3335 & ~n3898 ;
  assign n3900 = n3242 & ~n3890 ;
  assign n3901 = ~n3242 & ~n3894 ;
  assign n3902 = ~n3900 & ~n3901 ;
  assign n3903 = n3335 & ~n3902 ;
  assign n3904 = ~n3899 & ~n3903 ;
  assign n3905 = n3484 & ~n3904 ;
  assign n3906 = n3335 & ~n3898 ;
  assign n3907 = ~n3335 & ~n3902 ;
  assign n3908 = ~n3906 & ~n3907 ;
  assign n3909 = n3439 & ~n3908 ;
  assign n3910 = ~n3287 & ~n3896 ;
  assign n3911 = n3287 & ~n3886 ;
  assign n3912 = ~n3910 & ~n3911 ;
  assign n3913 = ~n3384 & ~n3912 ;
  assign n3914 = x4 & n3384 ;
  assign n3915 = ~n3913 & ~n3914 ;
  assign n3916 = ~n3439 & ~n3915 ;
  assign n3917 = ~n3909 & ~n3916 ;
  assign n3918 = ~n3484 & ~n3917 ;
  assign n3919 = ~n3905 & ~n3918 ;
  assign n3920 = x229 & ~n2640 ;
  assign n3921 = x197 & n2640 ;
  assign n3922 = ~n3920 & ~n3921 ;
  assign n3923 = n2693 & ~n3922 ;
  assign n3924 = x165 & ~n2693 ;
  assign n3925 = ~n3923 & ~n3924 ;
  assign n3926 = n2742 & ~n3925 ;
  assign n3927 = x197 & ~n2640 ;
  assign n3928 = x229 & n2640 ;
  assign n3929 = ~n3927 & ~n3928 ;
  assign n3930 = ~n2742 & ~n3929 ;
  assign n3931 = ~n3926 & ~n3930 ;
  assign n3932 = ~n2841 & ~n3931 ;
  assign n3933 = ~n2693 & ~n3922 ;
  assign n3934 = x165 & n2693 ;
  assign n3935 = ~n3933 & ~n3934 ;
  assign n3936 = ~n2791 & ~n3935 ;
  assign n3937 = x133 & n2791 ;
  assign n3938 = ~n3936 & ~n3937 ;
  assign n3939 = n2841 & ~n3938 ;
  assign n3940 = ~n3932 & ~n3939 ;
  assign n3941 = ~n2887 & ~n3940 ;
  assign n3942 = x101 & n2887 ;
  assign n3943 = ~n3941 & ~n3942 ;
  assign n3944 = n2989 & ~n3943 ;
  assign n3945 = n2841 & ~n3931 ;
  assign n3946 = ~n2841 & ~n3938 ;
  assign n3947 = ~n3945 & ~n3946 ;
  assign n3948 = n2944 & ~n3947 ;
  assign n3949 = n2742 & ~n3929 ;
  assign n3950 = ~n2742 & ~n3925 ;
  assign n3951 = ~n3949 & ~n3950 ;
  assign n3952 = ~n2944 & ~n3951 ;
  assign n3953 = ~n3948 & ~n3952 ;
  assign n3954 = ~n2989 & ~n3953 ;
  assign n3955 = ~n3944 & ~n3954 ;
  assign n3956 = ~n3035 & ~n3955 ;
  assign n3957 = x69 & n3035 ;
  assign n3958 = ~n3956 & ~n3957 ;
  assign n3959 = n3139 & ~n3958 ;
  assign n3960 = n2944 & ~n3951 ;
  assign n3961 = ~n2944 & ~n3947 ;
  assign n3962 = ~n3960 & ~n3961 ;
  assign n3963 = ~n3093 & ~n3962 ;
  assign n3964 = n2989 & ~n3953 ;
  assign n3965 = ~n2989 & ~n3943 ;
  assign n3966 = ~n3964 & ~n3965 ;
  assign n3967 = n3093 & ~n3966 ;
  assign n3968 = ~n3963 & ~n3967 ;
  assign n3969 = ~n3139 & ~n3968 ;
  assign n3970 = ~n3959 & ~n3969 ;
  assign n3971 = ~n3185 & ~n3970 ;
  assign n3972 = x37 & n3185 ;
  assign n3973 = ~n3971 & ~n3972 ;
  assign n3974 = ~n3287 & ~n3973 ;
  assign n3975 = n3093 & ~n3962 ;
  assign n3976 = ~n3093 & ~n3966 ;
  assign n3977 = ~n3975 & ~n3976 ;
  assign n3978 = ~n3242 & ~n3977 ;
  assign n3979 = n3139 & ~n3968 ;
  assign n3980 = ~n3139 & ~n3958 ;
  assign n3981 = ~n3979 & ~n3980 ;
  assign n3982 = n3242 & ~n3981 ;
  assign n3983 = ~n3978 & ~n3982 ;
  assign n3984 = n3287 & ~n3983 ;
  assign n3985 = ~n3974 & ~n3984 ;
  assign n3986 = ~n3335 & ~n3985 ;
  assign n3987 = n3242 & ~n3977 ;
  assign n3988 = ~n3242 & ~n3981 ;
  assign n3989 = ~n3987 & ~n3988 ;
  assign n3990 = n3335 & ~n3989 ;
  assign n3991 = ~n3986 & ~n3990 ;
  assign n3992 = n3484 & ~n3991 ;
  assign n3993 = n3335 & ~n3985 ;
  assign n3994 = ~n3335 & ~n3989 ;
  assign n3995 = ~n3993 & ~n3994 ;
  assign n3996 = n3439 & ~n3995 ;
  assign n3997 = ~n3287 & ~n3983 ;
  assign n3998 = n3287 & ~n3973 ;
  assign n3999 = ~n3997 & ~n3998 ;
  assign n4000 = ~n3384 & ~n3999 ;
  assign n4001 = x5 & n3384 ;
  assign n4002 = ~n4000 & ~n4001 ;
  assign n4003 = ~n3439 & ~n4002 ;
  assign n4004 = ~n3996 & ~n4003 ;
  assign n4005 = ~n3484 & ~n4004 ;
  assign n4006 = ~n3992 & ~n4005 ;
  assign n4007 = x230 & ~n2640 ;
  assign n4008 = x198 & n2640 ;
  assign n4009 = ~n4007 & ~n4008 ;
  assign n4010 = n2693 & ~n4009 ;
  assign n4011 = x166 & ~n2693 ;
  assign n4012 = ~n4010 & ~n4011 ;
  assign n4013 = n2742 & ~n4012 ;
  assign n4014 = x198 & ~n2640 ;
  assign n4015 = x230 & n2640 ;
  assign n4016 = ~n4014 & ~n4015 ;
  assign n4017 = ~n2742 & ~n4016 ;
  assign n4018 = ~n4013 & ~n4017 ;
  assign n4019 = ~n2841 & ~n4018 ;
  assign n4020 = ~n2693 & ~n4009 ;
  assign n4021 = x166 & n2693 ;
  assign n4022 = ~n4020 & ~n4021 ;
  assign n4023 = ~n2791 & ~n4022 ;
  assign n4024 = x134 & n2791 ;
  assign n4025 = ~n4023 & ~n4024 ;
  assign n4026 = n2841 & ~n4025 ;
  assign n4027 = ~n4019 & ~n4026 ;
  assign n4028 = ~n2887 & ~n4027 ;
  assign n4029 = x102 & n2887 ;
  assign n4030 = ~n4028 & ~n4029 ;
  assign n4031 = n2989 & ~n4030 ;
  assign n4032 = n2841 & ~n4018 ;
  assign n4033 = ~n2841 & ~n4025 ;
  assign n4034 = ~n4032 & ~n4033 ;
  assign n4035 = n2944 & ~n4034 ;
  assign n4036 = n2742 & ~n4016 ;
  assign n4037 = ~n2742 & ~n4012 ;
  assign n4038 = ~n4036 & ~n4037 ;
  assign n4039 = ~n2944 & ~n4038 ;
  assign n4040 = ~n4035 & ~n4039 ;
  assign n4041 = ~n2989 & ~n4040 ;
  assign n4042 = ~n4031 & ~n4041 ;
  assign n4043 = ~n3035 & ~n4042 ;
  assign n4044 = x70 & n3035 ;
  assign n4045 = ~n4043 & ~n4044 ;
  assign n4046 = n3139 & ~n4045 ;
  assign n4047 = n2944 & ~n4038 ;
  assign n4048 = ~n2944 & ~n4034 ;
  assign n4049 = ~n4047 & ~n4048 ;
  assign n4050 = ~n3093 & ~n4049 ;
  assign n4051 = n2989 & ~n4040 ;
  assign n4052 = ~n2989 & ~n4030 ;
  assign n4053 = ~n4051 & ~n4052 ;
  assign n4054 = n3093 & ~n4053 ;
  assign n4055 = ~n4050 & ~n4054 ;
  assign n4056 = ~n3139 & ~n4055 ;
  assign n4057 = ~n4046 & ~n4056 ;
  assign n4058 = ~n3185 & ~n4057 ;
  assign n4059 = x38 & n3185 ;
  assign n4060 = ~n4058 & ~n4059 ;
  assign n4061 = ~n3287 & ~n4060 ;
  assign n4062 = n3093 & ~n4049 ;
  assign n4063 = ~n3093 & ~n4053 ;
  assign n4064 = ~n4062 & ~n4063 ;
  assign n4065 = ~n3242 & ~n4064 ;
  assign n4066 = n3139 & ~n4055 ;
  assign n4067 = ~n3139 & ~n4045 ;
  assign n4068 = ~n4066 & ~n4067 ;
  assign n4069 = n3242 & ~n4068 ;
  assign n4070 = ~n4065 & ~n4069 ;
  assign n4071 = n3287 & ~n4070 ;
  assign n4072 = ~n4061 & ~n4071 ;
  assign n4073 = ~n3335 & ~n4072 ;
  assign n4074 = n3242 & ~n4064 ;
  assign n4075 = ~n3242 & ~n4068 ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = n3335 & ~n4076 ;
  assign n4078 = ~n4073 & ~n4077 ;
  assign n4079 = n3484 & ~n4078 ;
  assign n4080 = n3335 & ~n4072 ;
  assign n4081 = ~n3335 & ~n4076 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4083 = n3439 & ~n4082 ;
  assign n4084 = ~n3287 & ~n4070 ;
  assign n4085 = n3287 & ~n4060 ;
  assign n4086 = ~n4084 & ~n4085 ;
  assign n4087 = ~n3384 & ~n4086 ;
  assign n4088 = x6 & n3384 ;
  assign n4089 = ~n4087 & ~n4088 ;
  assign n4090 = ~n3439 & ~n4089 ;
  assign n4091 = ~n4083 & ~n4090 ;
  assign n4092 = ~n3484 & ~n4091 ;
  assign n4093 = ~n4079 & ~n4092 ;
  assign n4094 = x231 & ~n2640 ;
  assign n4095 = x199 & n2640 ;
  assign n4096 = ~n4094 & ~n4095 ;
  assign n4097 = n2693 & ~n4096 ;
  assign n4098 = x167 & ~n2693 ;
  assign n4099 = ~n4097 & ~n4098 ;
  assign n4100 = n2742 & ~n4099 ;
  assign n4101 = x199 & ~n2640 ;
  assign n4102 = x231 & n2640 ;
  assign n4103 = ~n4101 & ~n4102 ;
  assign n4104 = ~n2742 & ~n4103 ;
  assign n4105 = ~n4100 & ~n4104 ;
  assign n4106 = ~n2841 & ~n4105 ;
  assign n4107 = ~n2693 & ~n4096 ;
  assign n4108 = x167 & n2693 ;
  assign n4109 = ~n4107 & ~n4108 ;
  assign n4110 = ~n2791 & ~n4109 ;
  assign n4111 = x135 & n2791 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = n2841 & ~n4112 ;
  assign n4114 = ~n4106 & ~n4113 ;
  assign n4115 = ~n2887 & ~n4114 ;
  assign n4116 = x103 & n2887 ;
  assign n4117 = ~n4115 & ~n4116 ;
  assign n4118 = n2989 & ~n4117 ;
  assign n4119 = n2841 & ~n4105 ;
  assign n4120 = ~n2841 & ~n4112 ;
  assign n4121 = ~n4119 & ~n4120 ;
  assign n4122 = n2944 & ~n4121 ;
  assign n4123 = n2742 & ~n4103 ;
  assign n4124 = ~n2742 & ~n4099 ;
  assign n4125 = ~n4123 & ~n4124 ;
  assign n4126 = ~n2944 & ~n4125 ;
  assign n4127 = ~n4122 & ~n4126 ;
  assign n4128 = ~n2989 & ~n4127 ;
  assign n4129 = ~n4118 & ~n4128 ;
  assign n4130 = ~n3035 & ~n4129 ;
  assign n4131 = x71 & n3035 ;
  assign n4132 = ~n4130 & ~n4131 ;
  assign n4133 = n3139 & ~n4132 ;
  assign n4134 = n2944 & ~n4125 ;
  assign n4135 = ~n2944 & ~n4121 ;
  assign n4136 = ~n4134 & ~n4135 ;
  assign n4137 = ~n3093 & ~n4136 ;
  assign n4138 = n2989 & ~n4127 ;
  assign n4139 = ~n2989 & ~n4117 ;
  assign n4140 = ~n4138 & ~n4139 ;
  assign n4141 = n3093 & ~n4140 ;
  assign n4142 = ~n4137 & ~n4141 ;
  assign n4143 = ~n3139 & ~n4142 ;
  assign n4144 = ~n4133 & ~n4143 ;
  assign n4145 = ~n3185 & ~n4144 ;
  assign n4146 = x39 & n3185 ;
  assign n4147 = ~n4145 & ~n4146 ;
  assign n4148 = ~n3287 & ~n4147 ;
  assign n4149 = n3093 & ~n4136 ;
  assign n4150 = ~n3093 & ~n4140 ;
  assign n4151 = ~n4149 & ~n4150 ;
  assign n4152 = ~n3242 & ~n4151 ;
  assign n4153 = n3139 & ~n4142 ;
  assign n4154 = ~n3139 & ~n4132 ;
  assign n4155 = ~n4153 & ~n4154 ;
  assign n4156 = n3242 & ~n4155 ;
  assign n4157 = ~n4152 & ~n4156 ;
  assign n4158 = n3287 & ~n4157 ;
  assign n4159 = ~n4148 & ~n4158 ;
  assign n4160 = ~n3335 & ~n4159 ;
  assign n4161 = n3242 & ~n4151 ;
  assign n4162 = ~n3242 & ~n4155 ;
  assign n4163 = ~n4161 & ~n4162 ;
  assign n4164 = n3335 & ~n4163 ;
  assign n4165 = ~n4160 & ~n4164 ;
  assign n4166 = n3484 & ~n4165 ;
  assign n4167 = n3335 & ~n4159 ;
  assign n4168 = ~n3335 & ~n4163 ;
  assign n4169 = ~n4167 & ~n4168 ;
  assign n4170 = n3439 & ~n4169 ;
  assign n4171 = ~n3287 & ~n4157 ;
  assign n4172 = n3287 & ~n4147 ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4174 = ~n3384 & ~n4173 ;
  assign n4175 = x7 & n3384 ;
  assign n4176 = ~n4174 & ~n4175 ;
  assign n4177 = ~n3439 & ~n4176 ;
  assign n4178 = ~n4170 & ~n4177 ;
  assign n4179 = ~n3484 & ~n4178 ;
  assign n4180 = ~n4166 & ~n4179 ;
  assign n4181 = x232 & ~n2640 ;
  assign n4182 = x200 & n2640 ;
  assign n4183 = ~n4181 & ~n4182 ;
  assign n4184 = n2693 & ~n4183 ;
  assign n4185 = x168 & ~n2693 ;
  assign n4186 = ~n4184 & ~n4185 ;
  assign n4187 = n2742 & ~n4186 ;
  assign n4188 = x200 & ~n2640 ;
  assign n4189 = x232 & n2640 ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = ~n2742 & ~n4190 ;
  assign n4192 = ~n4187 & ~n4191 ;
  assign n4193 = ~n2841 & ~n4192 ;
  assign n4194 = ~n2693 & ~n4183 ;
  assign n4195 = x168 & n2693 ;
  assign n4196 = ~n4194 & ~n4195 ;
  assign n4197 = ~n2791 & ~n4196 ;
  assign n4198 = x136 & n2791 ;
  assign n4199 = ~n4197 & ~n4198 ;
  assign n4200 = n2841 & ~n4199 ;
  assign n4201 = ~n4193 & ~n4200 ;
  assign n4202 = ~n2887 & ~n4201 ;
  assign n4203 = x104 & n2887 ;
  assign n4204 = ~n4202 & ~n4203 ;
  assign n4205 = n2989 & ~n4204 ;
  assign n4206 = n2841 & ~n4192 ;
  assign n4207 = ~n2841 & ~n4199 ;
  assign n4208 = ~n4206 & ~n4207 ;
  assign n4209 = n2944 & ~n4208 ;
  assign n4210 = n2742 & ~n4190 ;
  assign n4211 = ~n2742 & ~n4186 ;
  assign n4212 = ~n4210 & ~n4211 ;
  assign n4213 = ~n2944 & ~n4212 ;
  assign n4214 = ~n4209 & ~n4213 ;
  assign n4215 = ~n2989 & ~n4214 ;
  assign n4216 = ~n4205 & ~n4215 ;
  assign n4217 = ~n3035 & ~n4216 ;
  assign n4218 = x72 & n3035 ;
  assign n4219 = ~n4217 & ~n4218 ;
  assign n4220 = n3139 & ~n4219 ;
  assign n4221 = n2944 & ~n4212 ;
  assign n4222 = ~n2944 & ~n4208 ;
  assign n4223 = ~n4221 & ~n4222 ;
  assign n4224 = ~n3093 & ~n4223 ;
  assign n4225 = n2989 & ~n4214 ;
  assign n4226 = ~n2989 & ~n4204 ;
  assign n4227 = ~n4225 & ~n4226 ;
  assign n4228 = n3093 & ~n4227 ;
  assign n4229 = ~n4224 & ~n4228 ;
  assign n4230 = ~n3139 & ~n4229 ;
  assign n4231 = ~n4220 & ~n4230 ;
  assign n4232 = ~n3185 & ~n4231 ;
  assign n4233 = x40 & n3185 ;
  assign n4234 = ~n4232 & ~n4233 ;
  assign n4235 = ~n3287 & ~n4234 ;
  assign n4236 = n3093 & ~n4223 ;
  assign n4237 = ~n3093 & ~n4227 ;
  assign n4238 = ~n4236 & ~n4237 ;
  assign n4239 = ~n3242 & ~n4238 ;
  assign n4240 = n3139 & ~n4229 ;
  assign n4241 = ~n3139 & ~n4219 ;
  assign n4242 = ~n4240 & ~n4241 ;
  assign n4243 = n3242 & ~n4242 ;
  assign n4244 = ~n4239 & ~n4243 ;
  assign n4245 = n3287 & ~n4244 ;
  assign n4246 = ~n4235 & ~n4245 ;
  assign n4247 = ~n3335 & ~n4246 ;
  assign n4248 = n3242 & ~n4238 ;
  assign n4249 = ~n3242 & ~n4242 ;
  assign n4250 = ~n4248 & ~n4249 ;
  assign n4251 = n3335 & ~n4250 ;
  assign n4252 = ~n4247 & ~n4251 ;
  assign n4253 = n3484 & ~n4252 ;
  assign n4254 = n3335 & ~n4246 ;
  assign n4255 = ~n3335 & ~n4250 ;
  assign n4256 = ~n4254 & ~n4255 ;
  assign n4257 = n3439 & ~n4256 ;
  assign n4258 = ~n3287 & ~n4244 ;
  assign n4259 = n3287 & ~n4234 ;
  assign n4260 = ~n4258 & ~n4259 ;
  assign n4261 = ~n3384 & ~n4260 ;
  assign n4262 = x8 & n3384 ;
  assign n4263 = ~n4261 & ~n4262 ;
  assign n4264 = ~n3439 & ~n4263 ;
  assign n4265 = ~n4257 & ~n4264 ;
  assign n4266 = ~n3484 & ~n4265 ;
  assign n4267 = ~n4253 & ~n4266 ;
  assign n4268 = x233 & ~n2640 ;
  assign n4269 = x201 & n2640 ;
  assign n4270 = ~n4268 & ~n4269 ;
  assign n4271 = n2693 & ~n4270 ;
  assign n4272 = x169 & ~n2693 ;
  assign n4273 = ~n4271 & ~n4272 ;
  assign n4274 = n2742 & ~n4273 ;
  assign n4275 = x201 & ~n2640 ;
  assign n4276 = x233 & n2640 ;
  assign n4277 = ~n4275 & ~n4276 ;
  assign n4278 = ~n2742 & ~n4277 ;
  assign n4279 = ~n4274 & ~n4278 ;
  assign n4280 = ~n2841 & ~n4279 ;
  assign n4281 = ~n2693 & ~n4270 ;
  assign n4282 = x169 & n2693 ;
  assign n4283 = ~n4281 & ~n4282 ;
  assign n4284 = ~n2791 & ~n4283 ;
  assign n4285 = x137 & n2791 ;
  assign n4286 = ~n4284 & ~n4285 ;
  assign n4287 = n2841 & ~n4286 ;
  assign n4288 = ~n4280 & ~n4287 ;
  assign n4289 = ~n2887 & ~n4288 ;
  assign n4290 = x105 & n2887 ;
  assign n4291 = ~n4289 & ~n4290 ;
  assign n4292 = n2989 & ~n4291 ;
  assign n4293 = n2841 & ~n4279 ;
  assign n4294 = ~n2841 & ~n4286 ;
  assign n4295 = ~n4293 & ~n4294 ;
  assign n4296 = n2944 & ~n4295 ;
  assign n4297 = n2742 & ~n4277 ;
  assign n4298 = ~n2742 & ~n4273 ;
  assign n4299 = ~n4297 & ~n4298 ;
  assign n4300 = ~n2944 & ~n4299 ;
  assign n4301 = ~n4296 & ~n4300 ;
  assign n4302 = ~n2989 & ~n4301 ;
  assign n4303 = ~n4292 & ~n4302 ;
  assign n4304 = ~n3035 & ~n4303 ;
  assign n4305 = x73 & n3035 ;
  assign n4306 = ~n4304 & ~n4305 ;
  assign n4307 = n3139 & ~n4306 ;
  assign n4308 = n2944 & ~n4299 ;
  assign n4309 = ~n2944 & ~n4295 ;
  assign n4310 = ~n4308 & ~n4309 ;
  assign n4311 = ~n3093 & ~n4310 ;
  assign n4312 = n2989 & ~n4301 ;
  assign n4313 = ~n2989 & ~n4291 ;
  assign n4314 = ~n4312 & ~n4313 ;
  assign n4315 = n3093 & ~n4314 ;
  assign n4316 = ~n4311 & ~n4315 ;
  assign n4317 = ~n3139 & ~n4316 ;
  assign n4318 = ~n4307 & ~n4317 ;
  assign n4319 = ~n3185 & ~n4318 ;
  assign n4320 = x41 & n3185 ;
  assign n4321 = ~n4319 & ~n4320 ;
  assign n4322 = ~n3287 & ~n4321 ;
  assign n4323 = n3093 & ~n4310 ;
  assign n4324 = ~n3093 & ~n4314 ;
  assign n4325 = ~n4323 & ~n4324 ;
  assign n4326 = ~n3242 & ~n4325 ;
  assign n4327 = n3139 & ~n4316 ;
  assign n4328 = ~n3139 & ~n4306 ;
  assign n4329 = ~n4327 & ~n4328 ;
  assign n4330 = n3242 & ~n4329 ;
  assign n4331 = ~n4326 & ~n4330 ;
  assign n4332 = n3287 & ~n4331 ;
  assign n4333 = ~n4322 & ~n4332 ;
  assign n4334 = ~n3335 & ~n4333 ;
  assign n4335 = n3242 & ~n4325 ;
  assign n4336 = ~n3242 & ~n4329 ;
  assign n4337 = ~n4335 & ~n4336 ;
  assign n4338 = n3335 & ~n4337 ;
  assign n4339 = ~n4334 & ~n4338 ;
  assign n4340 = n3484 & ~n4339 ;
  assign n4341 = n3335 & ~n4333 ;
  assign n4342 = ~n3335 & ~n4337 ;
  assign n4343 = ~n4341 & ~n4342 ;
  assign n4344 = n3439 & ~n4343 ;
  assign n4345 = ~n3287 & ~n4331 ;
  assign n4346 = n3287 & ~n4321 ;
  assign n4347 = ~n4345 & ~n4346 ;
  assign n4348 = ~n3384 & ~n4347 ;
  assign n4349 = x9 & n3384 ;
  assign n4350 = ~n4348 & ~n4349 ;
  assign n4351 = ~n3439 & ~n4350 ;
  assign n4352 = ~n4344 & ~n4351 ;
  assign n4353 = ~n3484 & ~n4352 ;
  assign n4354 = ~n4340 & ~n4353 ;
  assign n4355 = x234 & ~n2640 ;
  assign n4356 = x202 & n2640 ;
  assign n4357 = ~n4355 & ~n4356 ;
  assign n4358 = n2693 & ~n4357 ;
  assign n4359 = x170 & ~n2693 ;
  assign n4360 = ~n4358 & ~n4359 ;
  assign n4361 = n2742 & ~n4360 ;
  assign n4362 = x202 & ~n2640 ;
  assign n4363 = x234 & n2640 ;
  assign n4364 = ~n4362 & ~n4363 ;
  assign n4365 = ~n2742 & ~n4364 ;
  assign n4366 = ~n4361 & ~n4365 ;
  assign n4367 = ~n2841 & ~n4366 ;
  assign n4368 = ~n2693 & ~n4357 ;
  assign n4369 = x170 & n2693 ;
  assign n4370 = ~n4368 & ~n4369 ;
  assign n4371 = ~n2791 & ~n4370 ;
  assign n4372 = x138 & n2791 ;
  assign n4373 = ~n4371 & ~n4372 ;
  assign n4374 = n2841 & ~n4373 ;
  assign n4375 = ~n4367 & ~n4374 ;
  assign n4376 = ~n2887 & ~n4375 ;
  assign n4377 = x106 & n2887 ;
  assign n4378 = ~n4376 & ~n4377 ;
  assign n4379 = n2989 & ~n4378 ;
  assign n4380 = n2841 & ~n4366 ;
  assign n4381 = ~n2841 & ~n4373 ;
  assign n4382 = ~n4380 & ~n4381 ;
  assign n4383 = n2944 & ~n4382 ;
  assign n4384 = n2742 & ~n4364 ;
  assign n4385 = ~n2742 & ~n4360 ;
  assign n4386 = ~n4384 & ~n4385 ;
  assign n4387 = ~n2944 & ~n4386 ;
  assign n4388 = ~n4383 & ~n4387 ;
  assign n4389 = ~n2989 & ~n4388 ;
  assign n4390 = ~n4379 & ~n4389 ;
  assign n4391 = ~n3035 & ~n4390 ;
  assign n4392 = x74 & n3035 ;
  assign n4393 = ~n4391 & ~n4392 ;
  assign n4394 = n3139 & ~n4393 ;
  assign n4395 = n2944 & ~n4386 ;
  assign n4396 = ~n2944 & ~n4382 ;
  assign n4397 = ~n4395 & ~n4396 ;
  assign n4398 = ~n3093 & ~n4397 ;
  assign n4399 = n2989 & ~n4388 ;
  assign n4400 = ~n2989 & ~n4378 ;
  assign n4401 = ~n4399 & ~n4400 ;
  assign n4402 = n3093 & ~n4401 ;
  assign n4403 = ~n4398 & ~n4402 ;
  assign n4404 = ~n3139 & ~n4403 ;
  assign n4405 = ~n4394 & ~n4404 ;
  assign n4406 = ~n3185 & ~n4405 ;
  assign n4407 = x42 & n3185 ;
  assign n4408 = ~n4406 & ~n4407 ;
  assign n4409 = ~n3287 & ~n4408 ;
  assign n4410 = n3093 & ~n4397 ;
  assign n4411 = ~n3093 & ~n4401 ;
  assign n4412 = ~n4410 & ~n4411 ;
  assign n4413 = ~n3242 & ~n4412 ;
  assign n4414 = n3139 & ~n4403 ;
  assign n4415 = ~n3139 & ~n4393 ;
  assign n4416 = ~n4414 & ~n4415 ;
  assign n4417 = n3242 & ~n4416 ;
  assign n4418 = ~n4413 & ~n4417 ;
  assign n4419 = n3287 & ~n4418 ;
  assign n4420 = ~n4409 & ~n4419 ;
  assign n4421 = ~n3335 & ~n4420 ;
  assign n4422 = n3242 & ~n4412 ;
  assign n4423 = ~n3242 & ~n4416 ;
  assign n4424 = ~n4422 & ~n4423 ;
  assign n4425 = n3335 & ~n4424 ;
  assign n4426 = ~n4421 & ~n4425 ;
  assign n4427 = n3484 & ~n4426 ;
  assign n4428 = n3335 & ~n4420 ;
  assign n4429 = ~n3335 & ~n4424 ;
  assign n4430 = ~n4428 & ~n4429 ;
  assign n4431 = n3439 & ~n4430 ;
  assign n4432 = ~n3287 & ~n4418 ;
  assign n4433 = n3287 & ~n4408 ;
  assign n4434 = ~n4432 & ~n4433 ;
  assign n4435 = ~n3384 & ~n4434 ;
  assign n4436 = x10 & n3384 ;
  assign n4437 = ~n4435 & ~n4436 ;
  assign n4438 = ~n3439 & ~n4437 ;
  assign n4439 = ~n4431 & ~n4438 ;
  assign n4440 = ~n3484 & ~n4439 ;
  assign n4441 = ~n4427 & ~n4440 ;
  assign n4442 = x235 & ~n2640 ;
  assign n4443 = x203 & n2640 ;
  assign n4444 = ~n4442 & ~n4443 ;
  assign n4445 = n2693 & ~n4444 ;
  assign n4446 = x171 & ~n2693 ;
  assign n4447 = ~n4445 & ~n4446 ;
  assign n4448 = n2742 & ~n4447 ;
  assign n4449 = x203 & ~n2640 ;
  assign n4450 = x235 & n2640 ;
  assign n4451 = ~n4449 & ~n4450 ;
  assign n4452 = ~n2742 & ~n4451 ;
  assign n4453 = ~n4448 & ~n4452 ;
  assign n4454 = ~n2841 & ~n4453 ;
  assign n4455 = ~n2693 & ~n4444 ;
  assign n4456 = x171 & n2693 ;
  assign n4457 = ~n4455 & ~n4456 ;
  assign n4458 = ~n2791 & ~n4457 ;
  assign n4459 = x139 & n2791 ;
  assign n4460 = ~n4458 & ~n4459 ;
  assign n4461 = n2841 & ~n4460 ;
  assign n4462 = ~n4454 & ~n4461 ;
  assign n4463 = ~n2887 & ~n4462 ;
  assign n4464 = x107 & n2887 ;
  assign n4465 = ~n4463 & ~n4464 ;
  assign n4466 = n2989 & ~n4465 ;
  assign n4467 = n2841 & ~n4453 ;
  assign n4468 = ~n2841 & ~n4460 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = n2944 & ~n4469 ;
  assign n4471 = n2742 & ~n4451 ;
  assign n4472 = ~n2742 & ~n4447 ;
  assign n4473 = ~n4471 & ~n4472 ;
  assign n4474 = ~n2944 & ~n4473 ;
  assign n4475 = ~n4470 & ~n4474 ;
  assign n4476 = ~n2989 & ~n4475 ;
  assign n4477 = ~n4466 & ~n4476 ;
  assign n4478 = ~n3035 & ~n4477 ;
  assign n4479 = x75 & n3035 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = n3139 & ~n4480 ;
  assign n4482 = n2944 & ~n4473 ;
  assign n4483 = ~n2944 & ~n4469 ;
  assign n4484 = ~n4482 & ~n4483 ;
  assign n4485 = ~n3093 & ~n4484 ;
  assign n4486 = n2989 & ~n4475 ;
  assign n4487 = ~n2989 & ~n4465 ;
  assign n4488 = ~n4486 & ~n4487 ;
  assign n4489 = n3093 & ~n4488 ;
  assign n4490 = ~n4485 & ~n4489 ;
  assign n4491 = ~n3139 & ~n4490 ;
  assign n4492 = ~n4481 & ~n4491 ;
  assign n4493 = ~n3185 & ~n4492 ;
  assign n4494 = x43 & n3185 ;
  assign n4495 = ~n4493 & ~n4494 ;
  assign n4496 = ~n3287 & ~n4495 ;
  assign n4497 = n3093 & ~n4484 ;
  assign n4498 = ~n3093 & ~n4488 ;
  assign n4499 = ~n4497 & ~n4498 ;
  assign n4500 = ~n3242 & ~n4499 ;
  assign n4501 = n3139 & ~n4490 ;
  assign n4502 = ~n3139 & ~n4480 ;
  assign n4503 = ~n4501 & ~n4502 ;
  assign n4504 = n3242 & ~n4503 ;
  assign n4505 = ~n4500 & ~n4504 ;
  assign n4506 = n3287 & ~n4505 ;
  assign n4507 = ~n4496 & ~n4506 ;
  assign n4508 = ~n3335 & ~n4507 ;
  assign n4509 = n3242 & ~n4499 ;
  assign n4510 = ~n3242 & ~n4503 ;
  assign n4511 = ~n4509 & ~n4510 ;
  assign n4512 = n3335 & ~n4511 ;
  assign n4513 = ~n4508 & ~n4512 ;
  assign n4514 = n3484 & ~n4513 ;
  assign n4515 = n3335 & ~n4507 ;
  assign n4516 = ~n3335 & ~n4511 ;
  assign n4517 = ~n4515 & ~n4516 ;
  assign n4518 = n3439 & ~n4517 ;
  assign n4519 = ~n3287 & ~n4505 ;
  assign n4520 = n3287 & ~n4495 ;
  assign n4521 = ~n4519 & ~n4520 ;
  assign n4522 = ~n3384 & ~n4521 ;
  assign n4523 = x11 & n3384 ;
  assign n4524 = ~n4522 & ~n4523 ;
  assign n4525 = ~n3439 & ~n4524 ;
  assign n4526 = ~n4518 & ~n4525 ;
  assign n4527 = ~n3484 & ~n4526 ;
  assign n4528 = ~n4514 & ~n4527 ;
  assign n4529 = x236 & ~n2640 ;
  assign n4530 = x204 & n2640 ;
  assign n4531 = ~n4529 & ~n4530 ;
  assign n4532 = n2693 & ~n4531 ;
  assign n4533 = x172 & ~n2693 ;
  assign n4534 = ~n4532 & ~n4533 ;
  assign n4535 = n2742 & ~n4534 ;
  assign n4536 = x204 & ~n2640 ;
  assign n4537 = x236 & n2640 ;
  assign n4538 = ~n4536 & ~n4537 ;
  assign n4539 = ~n2742 & ~n4538 ;
  assign n4540 = ~n4535 & ~n4539 ;
  assign n4541 = ~n2841 & ~n4540 ;
  assign n4542 = ~n2693 & ~n4531 ;
  assign n4543 = x172 & n2693 ;
  assign n4544 = ~n4542 & ~n4543 ;
  assign n4545 = ~n2791 & ~n4544 ;
  assign n4546 = x140 & n2791 ;
  assign n4547 = ~n4545 & ~n4546 ;
  assign n4548 = n2841 & ~n4547 ;
  assign n4549 = ~n4541 & ~n4548 ;
  assign n4550 = ~n2887 & ~n4549 ;
  assign n4551 = x108 & n2887 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = n2989 & ~n4552 ;
  assign n4554 = n2841 & ~n4540 ;
  assign n4555 = ~n2841 & ~n4547 ;
  assign n4556 = ~n4554 & ~n4555 ;
  assign n4557 = n2944 & ~n4556 ;
  assign n4558 = n2742 & ~n4538 ;
  assign n4559 = ~n2742 & ~n4534 ;
  assign n4560 = ~n4558 & ~n4559 ;
  assign n4561 = ~n2944 & ~n4560 ;
  assign n4562 = ~n4557 & ~n4561 ;
  assign n4563 = ~n2989 & ~n4562 ;
  assign n4564 = ~n4553 & ~n4563 ;
  assign n4565 = ~n3035 & ~n4564 ;
  assign n4566 = x76 & n3035 ;
  assign n4567 = ~n4565 & ~n4566 ;
  assign n4568 = n3139 & ~n4567 ;
  assign n4569 = n2944 & ~n4560 ;
  assign n4570 = ~n2944 & ~n4556 ;
  assign n4571 = ~n4569 & ~n4570 ;
  assign n4572 = ~n3093 & ~n4571 ;
  assign n4573 = n2989 & ~n4562 ;
  assign n4574 = ~n2989 & ~n4552 ;
  assign n4575 = ~n4573 & ~n4574 ;
  assign n4576 = n3093 & ~n4575 ;
  assign n4577 = ~n4572 & ~n4576 ;
  assign n4578 = ~n3139 & ~n4577 ;
  assign n4579 = ~n4568 & ~n4578 ;
  assign n4580 = ~n3185 & ~n4579 ;
  assign n4581 = x44 & n3185 ;
  assign n4582 = ~n4580 & ~n4581 ;
  assign n4583 = ~n3287 & ~n4582 ;
  assign n4584 = n3093 & ~n4571 ;
  assign n4585 = ~n3093 & ~n4575 ;
  assign n4586 = ~n4584 & ~n4585 ;
  assign n4587 = ~n3242 & ~n4586 ;
  assign n4588 = n3139 & ~n4577 ;
  assign n4589 = ~n3139 & ~n4567 ;
  assign n4590 = ~n4588 & ~n4589 ;
  assign n4591 = n3242 & ~n4590 ;
  assign n4592 = ~n4587 & ~n4591 ;
  assign n4593 = n3287 & ~n4592 ;
  assign n4594 = ~n4583 & ~n4593 ;
  assign n4595 = ~n3335 & ~n4594 ;
  assign n4596 = n3242 & ~n4586 ;
  assign n4597 = ~n3242 & ~n4590 ;
  assign n4598 = ~n4596 & ~n4597 ;
  assign n4599 = n3335 & ~n4598 ;
  assign n4600 = ~n4595 & ~n4599 ;
  assign n4601 = n3484 & ~n4600 ;
  assign n4602 = n3335 & ~n4594 ;
  assign n4603 = ~n3335 & ~n4598 ;
  assign n4604 = ~n4602 & ~n4603 ;
  assign n4605 = n3439 & ~n4604 ;
  assign n4606 = ~n3287 & ~n4592 ;
  assign n4607 = n3287 & ~n4582 ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = ~n3384 & ~n4608 ;
  assign n4610 = x12 & n3384 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = ~n3439 & ~n4611 ;
  assign n4613 = ~n4605 & ~n4612 ;
  assign n4614 = ~n3484 & ~n4613 ;
  assign n4615 = ~n4601 & ~n4614 ;
  assign n4616 = x237 & ~n2640 ;
  assign n4617 = x205 & n2640 ;
  assign n4618 = ~n4616 & ~n4617 ;
  assign n4619 = n2693 & ~n4618 ;
  assign n4620 = x173 & ~n2693 ;
  assign n4621 = ~n4619 & ~n4620 ;
  assign n4622 = n2742 & ~n4621 ;
  assign n4623 = x205 & ~n2640 ;
  assign n4624 = x237 & n2640 ;
  assign n4625 = ~n4623 & ~n4624 ;
  assign n4626 = ~n2742 & ~n4625 ;
  assign n4627 = ~n4622 & ~n4626 ;
  assign n4628 = ~n2841 & ~n4627 ;
  assign n4629 = ~n2693 & ~n4618 ;
  assign n4630 = x173 & n2693 ;
  assign n4631 = ~n4629 & ~n4630 ;
  assign n4632 = ~n2791 & ~n4631 ;
  assign n4633 = x141 & n2791 ;
  assign n4634 = ~n4632 & ~n4633 ;
  assign n4635 = n2841 & ~n4634 ;
  assign n4636 = ~n4628 & ~n4635 ;
  assign n4637 = ~n2887 & ~n4636 ;
  assign n4638 = x109 & n2887 ;
  assign n4639 = ~n4637 & ~n4638 ;
  assign n4640 = n2989 & ~n4639 ;
  assign n4641 = n2841 & ~n4627 ;
  assign n4642 = ~n2841 & ~n4634 ;
  assign n4643 = ~n4641 & ~n4642 ;
  assign n4644 = n2944 & ~n4643 ;
  assign n4645 = n2742 & ~n4625 ;
  assign n4646 = ~n2742 & ~n4621 ;
  assign n4647 = ~n4645 & ~n4646 ;
  assign n4648 = ~n2944 & ~n4647 ;
  assign n4649 = ~n4644 & ~n4648 ;
  assign n4650 = ~n2989 & ~n4649 ;
  assign n4651 = ~n4640 & ~n4650 ;
  assign n4652 = ~n3035 & ~n4651 ;
  assign n4653 = x77 & n3035 ;
  assign n4654 = ~n4652 & ~n4653 ;
  assign n4655 = n3139 & ~n4654 ;
  assign n4656 = n2944 & ~n4647 ;
  assign n4657 = ~n2944 & ~n4643 ;
  assign n4658 = ~n4656 & ~n4657 ;
  assign n4659 = ~n3093 & ~n4658 ;
  assign n4660 = n2989 & ~n4649 ;
  assign n4661 = ~n2989 & ~n4639 ;
  assign n4662 = ~n4660 & ~n4661 ;
  assign n4663 = n3093 & ~n4662 ;
  assign n4664 = ~n4659 & ~n4663 ;
  assign n4665 = ~n3139 & ~n4664 ;
  assign n4666 = ~n4655 & ~n4665 ;
  assign n4667 = ~n3185 & ~n4666 ;
  assign n4668 = x45 & n3185 ;
  assign n4669 = ~n4667 & ~n4668 ;
  assign n4670 = ~n3287 & ~n4669 ;
  assign n4671 = n3093 & ~n4658 ;
  assign n4672 = ~n3093 & ~n4662 ;
  assign n4673 = ~n4671 & ~n4672 ;
  assign n4674 = ~n3242 & ~n4673 ;
  assign n4675 = n3139 & ~n4664 ;
  assign n4676 = ~n3139 & ~n4654 ;
  assign n4677 = ~n4675 & ~n4676 ;
  assign n4678 = n3242 & ~n4677 ;
  assign n4679 = ~n4674 & ~n4678 ;
  assign n4680 = n3287 & ~n4679 ;
  assign n4681 = ~n4670 & ~n4680 ;
  assign n4682 = ~n3335 & ~n4681 ;
  assign n4683 = n3242 & ~n4673 ;
  assign n4684 = ~n3242 & ~n4677 ;
  assign n4685 = ~n4683 & ~n4684 ;
  assign n4686 = n3335 & ~n4685 ;
  assign n4687 = ~n4682 & ~n4686 ;
  assign n4688 = n3484 & ~n4687 ;
  assign n4689 = n3335 & ~n4681 ;
  assign n4690 = ~n3335 & ~n4685 ;
  assign n4691 = ~n4689 & ~n4690 ;
  assign n4692 = n3439 & ~n4691 ;
  assign n4693 = ~n3287 & ~n4679 ;
  assign n4694 = n3287 & ~n4669 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = ~n3384 & ~n4695 ;
  assign n4697 = x13 & n3384 ;
  assign n4698 = ~n4696 & ~n4697 ;
  assign n4699 = ~n3439 & ~n4698 ;
  assign n4700 = ~n4692 & ~n4699 ;
  assign n4701 = ~n3484 & ~n4700 ;
  assign n4702 = ~n4688 & ~n4701 ;
  assign n4703 = x238 & ~n2640 ;
  assign n4704 = x206 & n2640 ;
  assign n4705 = ~n4703 & ~n4704 ;
  assign n4706 = n2693 & ~n4705 ;
  assign n4707 = x174 & ~n2693 ;
  assign n4708 = ~n4706 & ~n4707 ;
  assign n4709 = n2742 & ~n4708 ;
  assign n4710 = x206 & ~n2640 ;
  assign n4711 = x238 & n2640 ;
  assign n4712 = ~n4710 & ~n4711 ;
  assign n4713 = ~n2742 & ~n4712 ;
  assign n4714 = ~n4709 & ~n4713 ;
  assign n4715 = ~n2841 & ~n4714 ;
  assign n4716 = ~n2693 & ~n4705 ;
  assign n4717 = x174 & n2693 ;
  assign n4718 = ~n4716 & ~n4717 ;
  assign n4719 = ~n2791 & ~n4718 ;
  assign n4720 = x142 & n2791 ;
  assign n4721 = ~n4719 & ~n4720 ;
  assign n4722 = n2841 & ~n4721 ;
  assign n4723 = ~n4715 & ~n4722 ;
  assign n4724 = ~n2887 & ~n4723 ;
  assign n4725 = x110 & n2887 ;
  assign n4726 = ~n4724 & ~n4725 ;
  assign n4727 = n2989 & ~n4726 ;
  assign n4728 = n2841 & ~n4714 ;
  assign n4729 = ~n2841 & ~n4721 ;
  assign n4730 = ~n4728 & ~n4729 ;
  assign n4731 = n2944 & ~n4730 ;
  assign n4732 = n2742 & ~n4712 ;
  assign n4733 = ~n2742 & ~n4708 ;
  assign n4734 = ~n4732 & ~n4733 ;
  assign n4735 = ~n2944 & ~n4734 ;
  assign n4736 = ~n4731 & ~n4735 ;
  assign n4737 = ~n2989 & ~n4736 ;
  assign n4738 = ~n4727 & ~n4737 ;
  assign n4739 = ~n3035 & ~n4738 ;
  assign n4740 = x78 & n3035 ;
  assign n4741 = ~n4739 & ~n4740 ;
  assign n4742 = n3139 & ~n4741 ;
  assign n4743 = n2944 & ~n4734 ;
  assign n4744 = ~n2944 & ~n4730 ;
  assign n4745 = ~n4743 & ~n4744 ;
  assign n4746 = ~n3093 & ~n4745 ;
  assign n4747 = n2989 & ~n4736 ;
  assign n4748 = ~n2989 & ~n4726 ;
  assign n4749 = ~n4747 & ~n4748 ;
  assign n4750 = n3093 & ~n4749 ;
  assign n4751 = ~n4746 & ~n4750 ;
  assign n4752 = ~n3139 & ~n4751 ;
  assign n4753 = ~n4742 & ~n4752 ;
  assign n4754 = ~n3185 & ~n4753 ;
  assign n4755 = x46 & n3185 ;
  assign n4756 = ~n4754 & ~n4755 ;
  assign n4757 = ~n3287 & ~n4756 ;
  assign n4758 = n3093 & ~n4745 ;
  assign n4759 = ~n3093 & ~n4749 ;
  assign n4760 = ~n4758 & ~n4759 ;
  assign n4761 = ~n3242 & ~n4760 ;
  assign n4762 = n3139 & ~n4751 ;
  assign n4763 = ~n3139 & ~n4741 ;
  assign n4764 = ~n4762 & ~n4763 ;
  assign n4765 = n3242 & ~n4764 ;
  assign n4766 = ~n4761 & ~n4765 ;
  assign n4767 = n3287 & ~n4766 ;
  assign n4768 = ~n4757 & ~n4767 ;
  assign n4769 = ~n3335 & ~n4768 ;
  assign n4770 = n3242 & ~n4760 ;
  assign n4771 = ~n3242 & ~n4764 ;
  assign n4772 = ~n4770 & ~n4771 ;
  assign n4773 = n3335 & ~n4772 ;
  assign n4774 = ~n4769 & ~n4773 ;
  assign n4775 = n3484 & ~n4774 ;
  assign n4776 = n3335 & ~n4768 ;
  assign n4777 = ~n3335 & ~n4772 ;
  assign n4778 = ~n4776 & ~n4777 ;
  assign n4779 = n3439 & ~n4778 ;
  assign n4780 = ~n3287 & ~n4766 ;
  assign n4781 = n3287 & ~n4756 ;
  assign n4782 = ~n4780 & ~n4781 ;
  assign n4783 = ~n3384 & ~n4782 ;
  assign n4784 = x14 & n3384 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = ~n3439 & ~n4785 ;
  assign n4787 = ~n4779 & ~n4786 ;
  assign n4788 = ~n3484 & ~n4787 ;
  assign n4789 = ~n4775 & ~n4788 ;
  assign n4790 = x239 & ~n2640 ;
  assign n4791 = x207 & n2640 ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = n2693 & ~n4792 ;
  assign n4794 = x175 & ~n2693 ;
  assign n4795 = ~n4793 & ~n4794 ;
  assign n4796 = n2742 & ~n4795 ;
  assign n4797 = x207 & ~n2640 ;
  assign n4798 = x239 & n2640 ;
  assign n4799 = ~n4797 & ~n4798 ;
  assign n4800 = ~n2742 & ~n4799 ;
  assign n4801 = ~n4796 & ~n4800 ;
  assign n4802 = ~n2841 & ~n4801 ;
  assign n4803 = ~n2693 & ~n4792 ;
  assign n4804 = x175 & n2693 ;
  assign n4805 = ~n4803 & ~n4804 ;
  assign n4806 = ~n2791 & ~n4805 ;
  assign n4807 = x143 & n2791 ;
  assign n4808 = ~n4806 & ~n4807 ;
  assign n4809 = n2841 & ~n4808 ;
  assign n4810 = ~n4802 & ~n4809 ;
  assign n4811 = ~n2887 & ~n4810 ;
  assign n4812 = x111 & n2887 ;
  assign n4813 = ~n4811 & ~n4812 ;
  assign n4814 = n2989 & ~n4813 ;
  assign n4815 = n2841 & ~n4801 ;
  assign n4816 = ~n2841 & ~n4808 ;
  assign n4817 = ~n4815 & ~n4816 ;
  assign n4818 = n2944 & ~n4817 ;
  assign n4819 = n2742 & ~n4799 ;
  assign n4820 = ~n2742 & ~n4795 ;
  assign n4821 = ~n4819 & ~n4820 ;
  assign n4822 = ~n2944 & ~n4821 ;
  assign n4823 = ~n4818 & ~n4822 ;
  assign n4824 = ~n2989 & ~n4823 ;
  assign n4825 = ~n4814 & ~n4824 ;
  assign n4826 = ~n3035 & ~n4825 ;
  assign n4827 = x79 & n3035 ;
  assign n4828 = ~n4826 & ~n4827 ;
  assign n4829 = n3139 & ~n4828 ;
  assign n4830 = n2944 & ~n4821 ;
  assign n4831 = ~n2944 & ~n4817 ;
  assign n4832 = ~n4830 & ~n4831 ;
  assign n4833 = ~n3093 & ~n4832 ;
  assign n4834 = n2989 & ~n4823 ;
  assign n4835 = ~n2989 & ~n4813 ;
  assign n4836 = ~n4834 & ~n4835 ;
  assign n4837 = n3093 & ~n4836 ;
  assign n4838 = ~n4833 & ~n4837 ;
  assign n4839 = ~n3139 & ~n4838 ;
  assign n4840 = ~n4829 & ~n4839 ;
  assign n4841 = ~n3185 & ~n4840 ;
  assign n4842 = x47 & n3185 ;
  assign n4843 = ~n4841 & ~n4842 ;
  assign n4844 = ~n3287 & ~n4843 ;
  assign n4845 = n3093 & ~n4832 ;
  assign n4846 = ~n3093 & ~n4836 ;
  assign n4847 = ~n4845 & ~n4846 ;
  assign n4848 = ~n3242 & ~n4847 ;
  assign n4849 = n3139 & ~n4838 ;
  assign n4850 = ~n3139 & ~n4828 ;
  assign n4851 = ~n4849 & ~n4850 ;
  assign n4852 = n3242 & ~n4851 ;
  assign n4853 = ~n4848 & ~n4852 ;
  assign n4854 = n3287 & ~n4853 ;
  assign n4855 = ~n4844 & ~n4854 ;
  assign n4856 = ~n3335 & ~n4855 ;
  assign n4857 = n3242 & ~n4847 ;
  assign n4858 = ~n3242 & ~n4851 ;
  assign n4859 = ~n4857 & ~n4858 ;
  assign n4860 = n3335 & ~n4859 ;
  assign n4861 = ~n4856 & ~n4860 ;
  assign n4862 = n3484 & ~n4861 ;
  assign n4863 = n3335 & ~n4855 ;
  assign n4864 = ~n3335 & ~n4859 ;
  assign n4865 = ~n4863 & ~n4864 ;
  assign n4866 = n3439 & ~n4865 ;
  assign n4867 = ~n3287 & ~n4853 ;
  assign n4868 = n3287 & ~n4843 ;
  assign n4869 = ~n4867 & ~n4868 ;
  assign n4870 = ~n3384 & ~n4869 ;
  assign n4871 = x15 & n3384 ;
  assign n4872 = ~n4870 & ~n4871 ;
  assign n4873 = ~n3439 & ~n4872 ;
  assign n4874 = ~n4866 & ~n4873 ;
  assign n4875 = ~n3484 & ~n4874 ;
  assign n4876 = ~n4862 & ~n4875 ;
  assign n4877 = x240 & ~n2640 ;
  assign n4878 = x208 & n2640 ;
  assign n4879 = ~n4877 & ~n4878 ;
  assign n4880 = n2693 & ~n4879 ;
  assign n4881 = x176 & ~n2693 ;
  assign n4882 = ~n4880 & ~n4881 ;
  assign n4883 = n2742 & ~n4882 ;
  assign n4884 = x208 & ~n2640 ;
  assign n4885 = x240 & n2640 ;
  assign n4886 = ~n4884 & ~n4885 ;
  assign n4887 = ~n2742 & ~n4886 ;
  assign n4888 = ~n4883 & ~n4887 ;
  assign n4889 = ~n2841 & ~n4888 ;
  assign n4890 = ~n2693 & ~n4879 ;
  assign n4891 = x176 & n2693 ;
  assign n4892 = ~n4890 & ~n4891 ;
  assign n4893 = ~n2791 & ~n4892 ;
  assign n4894 = x144 & n2791 ;
  assign n4895 = ~n4893 & ~n4894 ;
  assign n4896 = n2841 & ~n4895 ;
  assign n4897 = ~n4889 & ~n4896 ;
  assign n4898 = ~n2887 & ~n4897 ;
  assign n4899 = x112 & n2887 ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = n2989 & ~n4900 ;
  assign n4902 = n2841 & ~n4888 ;
  assign n4903 = ~n2841 & ~n4895 ;
  assign n4904 = ~n4902 & ~n4903 ;
  assign n4905 = n2944 & ~n4904 ;
  assign n4906 = n2742 & ~n4886 ;
  assign n4907 = ~n2742 & ~n4882 ;
  assign n4908 = ~n4906 & ~n4907 ;
  assign n4909 = ~n2944 & ~n4908 ;
  assign n4910 = ~n4905 & ~n4909 ;
  assign n4911 = ~n2989 & ~n4910 ;
  assign n4912 = ~n4901 & ~n4911 ;
  assign n4913 = ~n3035 & ~n4912 ;
  assign n4914 = x80 & n3035 ;
  assign n4915 = ~n4913 & ~n4914 ;
  assign n4916 = n3139 & ~n4915 ;
  assign n4917 = n2944 & ~n4908 ;
  assign n4918 = ~n2944 & ~n4904 ;
  assign n4919 = ~n4917 & ~n4918 ;
  assign n4920 = ~n3093 & ~n4919 ;
  assign n4921 = n2989 & ~n4910 ;
  assign n4922 = ~n2989 & ~n4900 ;
  assign n4923 = ~n4921 & ~n4922 ;
  assign n4924 = n3093 & ~n4923 ;
  assign n4925 = ~n4920 & ~n4924 ;
  assign n4926 = ~n3139 & ~n4925 ;
  assign n4927 = ~n4916 & ~n4926 ;
  assign n4928 = ~n3185 & ~n4927 ;
  assign n4929 = x48 & n3185 ;
  assign n4930 = ~n4928 & ~n4929 ;
  assign n4931 = ~n3287 & ~n4930 ;
  assign n4932 = n3093 & ~n4919 ;
  assign n4933 = ~n3093 & ~n4923 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = ~n3242 & ~n4934 ;
  assign n4936 = n3139 & ~n4925 ;
  assign n4937 = ~n3139 & ~n4915 ;
  assign n4938 = ~n4936 & ~n4937 ;
  assign n4939 = n3242 & ~n4938 ;
  assign n4940 = ~n4935 & ~n4939 ;
  assign n4941 = n3287 & ~n4940 ;
  assign n4942 = ~n4931 & ~n4941 ;
  assign n4943 = ~n3335 & ~n4942 ;
  assign n4944 = n3242 & ~n4934 ;
  assign n4945 = ~n3242 & ~n4938 ;
  assign n4946 = ~n4944 & ~n4945 ;
  assign n4947 = n3335 & ~n4946 ;
  assign n4948 = ~n4943 & ~n4947 ;
  assign n4949 = n3484 & ~n4948 ;
  assign n4950 = n3335 & ~n4942 ;
  assign n4951 = ~n3335 & ~n4946 ;
  assign n4952 = ~n4950 & ~n4951 ;
  assign n4953 = n3439 & ~n4952 ;
  assign n4954 = ~n3287 & ~n4940 ;
  assign n4955 = n3287 & ~n4930 ;
  assign n4956 = ~n4954 & ~n4955 ;
  assign n4957 = ~n3384 & ~n4956 ;
  assign n4958 = x16 & n3384 ;
  assign n4959 = ~n4957 & ~n4958 ;
  assign n4960 = ~n3439 & ~n4959 ;
  assign n4961 = ~n4953 & ~n4960 ;
  assign n4962 = ~n3484 & ~n4961 ;
  assign n4963 = ~n4949 & ~n4962 ;
  assign n4964 = x241 & ~n2640 ;
  assign n4965 = x209 & n2640 ;
  assign n4966 = ~n4964 & ~n4965 ;
  assign n4967 = n2693 & ~n4966 ;
  assign n4968 = x177 & ~n2693 ;
  assign n4969 = ~n4967 & ~n4968 ;
  assign n4970 = n2742 & ~n4969 ;
  assign n4971 = x209 & ~n2640 ;
  assign n4972 = x241 & n2640 ;
  assign n4973 = ~n4971 & ~n4972 ;
  assign n4974 = ~n2742 & ~n4973 ;
  assign n4975 = ~n4970 & ~n4974 ;
  assign n4976 = ~n2841 & ~n4975 ;
  assign n4977 = ~n2693 & ~n4966 ;
  assign n4978 = x177 & n2693 ;
  assign n4979 = ~n4977 & ~n4978 ;
  assign n4980 = ~n2791 & ~n4979 ;
  assign n4981 = x145 & n2791 ;
  assign n4982 = ~n4980 & ~n4981 ;
  assign n4983 = n2841 & ~n4982 ;
  assign n4984 = ~n4976 & ~n4983 ;
  assign n4985 = ~n2887 & ~n4984 ;
  assign n4986 = x113 & n2887 ;
  assign n4987 = ~n4985 & ~n4986 ;
  assign n4988 = n2989 & ~n4987 ;
  assign n4989 = n2841 & ~n4975 ;
  assign n4990 = ~n2841 & ~n4982 ;
  assign n4991 = ~n4989 & ~n4990 ;
  assign n4992 = n2944 & ~n4991 ;
  assign n4993 = n2742 & ~n4973 ;
  assign n4994 = ~n2742 & ~n4969 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = ~n2944 & ~n4995 ;
  assign n4997 = ~n4992 & ~n4996 ;
  assign n4998 = ~n2989 & ~n4997 ;
  assign n4999 = ~n4988 & ~n4998 ;
  assign n5000 = ~n3035 & ~n4999 ;
  assign n5001 = x81 & n3035 ;
  assign n5002 = ~n5000 & ~n5001 ;
  assign n5003 = n3139 & ~n5002 ;
  assign n5004 = n2944 & ~n4995 ;
  assign n5005 = ~n2944 & ~n4991 ;
  assign n5006 = ~n5004 & ~n5005 ;
  assign n5007 = ~n3093 & ~n5006 ;
  assign n5008 = n2989 & ~n4997 ;
  assign n5009 = ~n2989 & ~n4987 ;
  assign n5010 = ~n5008 & ~n5009 ;
  assign n5011 = n3093 & ~n5010 ;
  assign n5012 = ~n5007 & ~n5011 ;
  assign n5013 = ~n3139 & ~n5012 ;
  assign n5014 = ~n5003 & ~n5013 ;
  assign n5015 = ~n3185 & ~n5014 ;
  assign n5016 = x49 & n3185 ;
  assign n5017 = ~n5015 & ~n5016 ;
  assign n5018 = ~n3287 & ~n5017 ;
  assign n5019 = n3093 & ~n5006 ;
  assign n5020 = ~n3093 & ~n5010 ;
  assign n5021 = ~n5019 & ~n5020 ;
  assign n5022 = ~n3242 & ~n5021 ;
  assign n5023 = n3139 & ~n5012 ;
  assign n5024 = ~n3139 & ~n5002 ;
  assign n5025 = ~n5023 & ~n5024 ;
  assign n5026 = n3242 & ~n5025 ;
  assign n5027 = ~n5022 & ~n5026 ;
  assign n5028 = n3287 & ~n5027 ;
  assign n5029 = ~n5018 & ~n5028 ;
  assign n5030 = ~n3335 & ~n5029 ;
  assign n5031 = n3242 & ~n5021 ;
  assign n5032 = ~n3242 & ~n5025 ;
  assign n5033 = ~n5031 & ~n5032 ;
  assign n5034 = n3335 & ~n5033 ;
  assign n5035 = ~n5030 & ~n5034 ;
  assign n5036 = n3484 & ~n5035 ;
  assign n5037 = n3335 & ~n5029 ;
  assign n5038 = ~n3335 & ~n5033 ;
  assign n5039 = ~n5037 & ~n5038 ;
  assign n5040 = n3439 & ~n5039 ;
  assign n5041 = ~n3287 & ~n5027 ;
  assign n5042 = n3287 & ~n5017 ;
  assign n5043 = ~n5041 & ~n5042 ;
  assign n5044 = ~n3384 & ~n5043 ;
  assign n5045 = x17 & n3384 ;
  assign n5046 = ~n5044 & ~n5045 ;
  assign n5047 = ~n3439 & ~n5046 ;
  assign n5048 = ~n5040 & ~n5047 ;
  assign n5049 = ~n3484 & ~n5048 ;
  assign n5050 = ~n5036 & ~n5049 ;
  assign n5051 = x242 & ~n2640 ;
  assign n5052 = x210 & n2640 ;
  assign n5053 = ~n5051 & ~n5052 ;
  assign n5054 = n2693 & ~n5053 ;
  assign n5055 = x178 & ~n2693 ;
  assign n5056 = ~n5054 & ~n5055 ;
  assign n5057 = n2742 & ~n5056 ;
  assign n5058 = x210 & ~n2640 ;
  assign n5059 = x242 & n2640 ;
  assign n5060 = ~n5058 & ~n5059 ;
  assign n5061 = ~n2742 & ~n5060 ;
  assign n5062 = ~n5057 & ~n5061 ;
  assign n5063 = ~n2841 & ~n5062 ;
  assign n5064 = ~n2693 & ~n5053 ;
  assign n5065 = x178 & n2693 ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = ~n2791 & ~n5066 ;
  assign n5068 = x146 & n2791 ;
  assign n5069 = ~n5067 & ~n5068 ;
  assign n5070 = n2841 & ~n5069 ;
  assign n5071 = ~n5063 & ~n5070 ;
  assign n5072 = ~n2887 & ~n5071 ;
  assign n5073 = x114 & n2887 ;
  assign n5074 = ~n5072 & ~n5073 ;
  assign n5075 = n2989 & ~n5074 ;
  assign n5076 = n2841 & ~n5062 ;
  assign n5077 = ~n2841 & ~n5069 ;
  assign n5078 = ~n5076 & ~n5077 ;
  assign n5079 = n2944 & ~n5078 ;
  assign n5080 = n2742 & ~n5060 ;
  assign n5081 = ~n2742 & ~n5056 ;
  assign n5082 = ~n5080 & ~n5081 ;
  assign n5083 = ~n2944 & ~n5082 ;
  assign n5084 = ~n5079 & ~n5083 ;
  assign n5085 = ~n2989 & ~n5084 ;
  assign n5086 = ~n5075 & ~n5085 ;
  assign n5087 = ~n3035 & ~n5086 ;
  assign n5088 = x82 & n3035 ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5090 = n3139 & ~n5089 ;
  assign n5091 = n2944 & ~n5082 ;
  assign n5092 = ~n2944 & ~n5078 ;
  assign n5093 = ~n5091 & ~n5092 ;
  assign n5094 = ~n3093 & ~n5093 ;
  assign n5095 = n2989 & ~n5084 ;
  assign n5096 = ~n2989 & ~n5074 ;
  assign n5097 = ~n5095 & ~n5096 ;
  assign n5098 = n3093 & ~n5097 ;
  assign n5099 = ~n5094 & ~n5098 ;
  assign n5100 = ~n3139 & ~n5099 ;
  assign n5101 = ~n5090 & ~n5100 ;
  assign n5102 = ~n3185 & ~n5101 ;
  assign n5103 = x50 & n3185 ;
  assign n5104 = ~n5102 & ~n5103 ;
  assign n5105 = ~n3287 & ~n5104 ;
  assign n5106 = n3093 & ~n5093 ;
  assign n5107 = ~n3093 & ~n5097 ;
  assign n5108 = ~n5106 & ~n5107 ;
  assign n5109 = ~n3242 & ~n5108 ;
  assign n5110 = n3139 & ~n5099 ;
  assign n5111 = ~n3139 & ~n5089 ;
  assign n5112 = ~n5110 & ~n5111 ;
  assign n5113 = n3242 & ~n5112 ;
  assign n5114 = ~n5109 & ~n5113 ;
  assign n5115 = n3287 & ~n5114 ;
  assign n5116 = ~n5105 & ~n5115 ;
  assign n5117 = ~n3335 & ~n5116 ;
  assign n5118 = n3242 & ~n5108 ;
  assign n5119 = ~n3242 & ~n5112 ;
  assign n5120 = ~n5118 & ~n5119 ;
  assign n5121 = n3335 & ~n5120 ;
  assign n5122 = ~n5117 & ~n5121 ;
  assign n5123 = n3484 & ~n5122 ;
  assign n5124 = n3335 & ~n5116 ;
  assign n5125 = ~n3335 & ~n5120 ;
  assign n5126 = ~n5124 & ~n5125 ;
  assign n5127 = n3439 & ~n5126 ;
  assign n5128 = ~n3287 & ~n5114 ;
  assign n5129 = n3287 & ~n5104 ;
  assign n5130 = ~n5128 & ~n5129 ;
  assign n5131 = ~n3384 & ~n5130 ;
  assign n5132 = x18 & n3384 ;
  assign n5133 = ~n5131 & ~n5132 ;
  assign n5134 = ~n3439 & ~n5133 ;
  assign n5135 = ~n5127 & ~n5134 ;
  assign n5136 = ~n3484 & ~n5135 ;
  assign n5137 = ~n5123 & ~n5136 ;
  assign n5138 = x243 & ~n2640 ;
  assign n5139 = x211 & n2640 ;
  assign n5140 = ~n5138 & ~n5139 ;
  assign n5141 = n2693 & ~n5140 ;
  assign n5142 = x179 & ~n2693 ;
  assign n5143 = ~n5141 & ~n5142 ;
  assign n5144 = n2742 & ~n5143 ;
  assign n5145 = x211 & ~n2640 ;
  assign n5146 = x243 & n2640 ;
  assign n5147 = ~n5145 & ~n5146 ;
  assign n5148 = ~n2742 & ~n5147 ;
  assign n5149 = ~n5144 & ~n5148 ;
  assign n5150 = ~n2841 & ~n5149 ;
  assign n5151 = ~n2693 & ~n5140 ;
  assign n5152 = x179 & n2693 ;
  assign n5153 = ~n5151 & ~n5152 ;
  assign n5154 = ~n2791 & ~n5153 ;
  assign n5155 = x147 & n2791 ;
  assign n5156 = ~n5154 & ~n5155 ;
  assign n5157 = n2841 & ~n5156 ;
  assign n5158 = ~n5150 & ~n5157 ;
  assign n5159 = ~n2887 & ~n5158 ;
  assign n5160 = x115 & n2887 ;
  assign n5161 = ~n5159 & ~n5160 ;
  assign n5162 = n2989 & ~n5161 ;
  assign n5163 = n2841 & ~n5149 ;
  assign n5164 = ~n2841 & ~n5156 ;
  assign n5165 = ~n5163 & ~n5164 ;
  assign n5166 = n2944 & ~n5165 ;
  assign n5167 = n2742 & ~n5147 ;
  assign n5168 = ~n2742 & ~n5143 ;
  assign n5169 = ~n5167 & ~n5168 ;
  assign n5170 = ~n2944 & ~n5169 ;
  assign n5171 = ~n5166 & ~n5170 ;
  assign n5172 = ~n2989 & ~n5171 ;
  assign n5173 = ~n5162 & ~n5172 ;
  assign n5174 = ~n3035 & ~n5173 ;
  assign n5175 = x83 & n3035 ;
  assign n5176 = ~n5174 & ~n5175 ;
  assign n5177 = n3139 & ~n5176 ;
  assign n5178 = n2944 & ~n5169 ;
  assign n5179 = ~n2944 & ~n5165 ;
  assign n5180 = ~n5178 & ~n5179 ;
  assign n5181 = ~n3093 & ~n5180 ;
  assign n5182 = n2989 & ~n5171 ;
  assign n5183 = ~n2989 & ~n5161 ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = n3093 & ~n5184 ;
  assign n5186 = ~n5181 & ~n5185 ;
  assign n5187 = ~n3139 & ~n5186 ;
  assign n5188 = ~n5177 & ~n5187 ;
  assign n5189 = ~n3185 & ~n5188 ;
  assign n5190 = x51 & n3185 ;
  assign n5191 = ~n5189 & ~n5190 ;
  assign n5192 = ~n3287 & ~n5191 ;
  assign n5193 = n3093 & ~n5180 ;
  assign n5194 = ~n3093 & ~n5184 ;
  assign n5195 = ~n5193 & ~n5194 ;
  assign n5196 = ~n3242 & ~n5195 ;
  assign n5197 = n3139 & ~n5186 ;
  assign n5198 = ~n3139 & ~n5176 ;
  assign n5199 = ~n5197 & ~n5198 ;
  assign n5200 = n3242 & ~n5199 ;
  assign n5201 = ~n5196 & ~n5200 ;
  assign n5202 = n3287 & ~n5201 ;
  assign n5203 = ~n5192 & ~n5202 ;
  assign n5204 = ~n3335 & ~n5203 ;
  assign n5205 = n3242 & ~n5195 ;
  assign n5206 = ~n3242 & ~n5199 ;
  assign n5207 = ~n5205 & ~n5206 ;
  assign n5208 = n3335 & ~n5207 ;
  assign n5209 = ~n5204 & ~n5208 ;
  assign n5210 = n3484 & ~n5209 ;
  assign n5211 = n3335 & ~n5203 ;
  assign n5212 = ~n3335 & ~n5207 ;
  assign n5213 = ~n5211 & ~n5212 ;
  assign n5214 = n3439 & ~n5213 ;
  assign n5215 = ~n3287 & ~n5201 ;
  assign n5216 = n3287 & ~n5191 ;
  assign n5217 = ~n5215 & ~n5216 ;
  assign n5218 = ~n3384 & ~n5217 ;
  assign n5219 = x19 & n3384 ;
  assign n5220 = ~n5218 & ~n5219 ;
  assign n5221 = ~n3439 & ~n5220 ;
  assign n5222 = ~n5214 & ~n5221 ;
  assign n5223 = ~n3484 & ~n5222 ;
  assign n5224 = ~n5210 & ~n5223 ;
  assign n5225 = x244 & ~n2640 ;
  assign n5226 = x212 & n2640 ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5228 = n2693 & ~n5227 ;
  assign n5229 = x180 & ~n2693 ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5231 = n2742 & ~n5230 ;
  assign n5232 = x212 & ~n2640 ;
  assign n5233 = x244 & n2640 ;
  assign n5234 = ~n5232 & ~n5233 ;
  assign n5235 = ~n2742 & ~n5234 ;
  assign n5236 = ~n5231 & ~n5235 ;
  assign n5237 = ~n2841 & ~n5236 ;
  assign n5238 = ~n2693 & ~n5227 ;
  assign n5239 = x180 & n2693 ;
  assign n5240 = ~n5238 & ~n5239 ;
  assign n5241 = ~n2791 & ~n5240 ;
  assign n5242 = x148 & n2791 ;
  assign n5243 = ~n5241 & ~n5242 ;
  assign n5244 = n2841 & ~n5243 ;
  assign n5245 = ~n5237 & ~n5244 ;
  assign n5246 = ~n2887 & ~n5245 ;
  assign n5247 = x116 & n2887 ;
  assign n5248 = ~n5246 & ~n5247 ;
  assign n5249 = n2989 & ~n5248 ;
  assign n5250 = n2841 & ~n5236 ;
  assign n5251 = ~n2841 & ~n5243 ;
  assign n5252 = ~n5250 & ~n5251 ;
  assign n5253 = n2944 & ~n5252 ;
  assign n5254 = n2742 & ~n5234 ;
  assign n5255 = ~n2742 & ~n5230 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = ~n2944 & ~n5256 ;
  assign n5258 = ~n5253 & ~n5257 ;
  assign n5259 = ~n2989 & ~n5258 ;
  assign n5260 = ~n5249 & ~n5259 ;
  assign n5261 = ~n3035 & ~n5260 ;
  assign n5262 = x84 & n3035 ;
  assign n5263 = ~n5261 & ~n5262 ;
  assign n5264 = n3139 & ~n5263 ;
  assign n5265 = n2944 & ~n5256 ;
  assign n5266 = ~n2944 & ~n5252 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = ~n3093 & ~n5267 ;
  assign n5269 = n2989 & ~n5258 ;
  assign n5270 = ~n2989 & ~n5248 ;
  assign n5271 = ~n5269 & ~n5270 ;
  assign n5272 = n3093 & ~n5271 ;
  assign n5273 = ~n5268 & ~n5272 ;
  assign n5274 = ~n3139 & ~n5273 ;
  assign n5275 = ~n5264 & ~n5274 ;
  assign n5276 = ~n3185 & ~n5275 ;
  assign n5277 = x52 & n3185 ;
  assign n5278 = ~n5276 & ~n5277 ;
  assign n5279 = ~n3287 & ~n5278 ;
  assign n5280 = n3093 & ~n5267 ;
  assign n5281 = ~n3093 & ~n5271 ;
  assign n5282 = ~n5280 & ~n5281 ;
  assign n5283 = ~n3242 & ~n5282 ;
  assign n5284 = n3139 & ~n5273 ;
  assign n5285 = ~n3139 & ~n5263 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = n3242 & ~n5286 ;
  assign n5288 = ~n5283 & ~n5287 ;
  assign n5289 = n3287 & ~n5288 ;
  assign n5290 = ~n5279 & ~n5289 ;
  assign n5291 = ~n3335 & ~n5290 ;
  assign n5292 = n3242 & ~n5282 ;
  assign n5293 = ~n3242 & ~n5286 ;
  assign n5294 = ~n5292 & ~n5293 ;
  assign n5295 = n3335 & ~n5294 ;
  assign n5296 = ~n5291 & ~n5295 ;
  assign n5297 = n3484 & ~n5296 ;
  assign n5298 = n3335 & ~n5290 ;
  assign n5299 = ~n3335 & ~n5294 ;
  assign n5300 = ~n5298 & ~n5299 ;
  assign n5301 = n3439 & ~n5300 ;
  assign n5302 = ~n3287 & ~n5288 ;
  assign n5303 = n3287 & ~n5278 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = ~n3384 & ~n5304 ;
  assign n5306 = x20 & n3384 ;
  assign n5307 = ~n5305 & ~n5306 ;
  assign n5308 = ~n3439 & ~n5307 ;
  assign n5309 = ~n5301 & ~n5308 ;
  assign n5310 = ~n3484 & ~n5309 ;
  assign n5311 = ~n5297 & ~n5310 ;
  assign n5312 = x245 & ~n2640 ;
  assign n5313 = x213 & n2640 ;
  assign n5314 = ~n5312 & ~n5313 ;
  assign n5315 = n2693 & ~n5314 ;
  assign n5316 = x181 & ~n2693 ;
  assign n5317 = ~n5315 & ~n5316 ;
  assign n5318 = n2742 & ~n5317 ;
  assign n5319 = x213 & ~n2640 ;
  assign n5320 = x245 & n2640 ;
  assign n5321 = ~n5319 & ~n5320 ;
  assign n5322 = ~n2742 & ~n5321 ;
  assign n5323 = ~n5318 & ~n5322 ;
  assign n5324 = ~n2841 & ~n5323 ;
  assign n5325 = ~n2693 & ~n5314 ;
  assign n5326 = x181 & n2693 ;
  assign n5327 = ~n5325 & ~n5326 ;
  assign n5328 = ~n2791 & ~n5327 ;
  assign n5329 = x149 & n2791 ;
  assign n5330 = ~n5328 & ~n5329 ;
  assign n5331 = n2841 & ~n5330 ;
  assign n5332 = ~n5324 & ~n5331 ;
  assign n5333 = ~n2887 & ~n5332 ;
  assign n5334 = x117 & n2887 ;
  assign n5335 = ~n5333 & ~n5334 ;
  assign n5336 = n2989 & ~n5335 ;
  assign n5337 = n2841 & ~n5323 ;
  assign n5338 = ~n2841 & ~n5330 ;
  assign n5339 = ~n5337 & ~n5338 ;
  assign n5340 = n2944 & ~n5339 ;
  assign n5341 = n2742 & ~n5321 ;
  assign n5342 = ~n2742 & ~n5317 ;
  assign n5343 = ~n5341 & ~n5342 ;
  assign n5344 = ~n2944 & ~n5343 ;
  assign n5345 = ~n5340 & ~n5344 ;
  assign n5346 = ~n2989 & ~n5345 ;
  assign n5347 = ~n5336 & ~n5346 ;
  assign n5348 = ~n3035 & ~n5347 ;
  assign n5349 = x85 & n3035 ;
  assign n5350 = ~n5348 & ~n5349 ;
  assign n5351 = n3139 & ~n5350 ;
  assign n5352 = n2944 & ~n5343 ;
  assign n5353 = ~n2944 & ~n5339 ;
  assign n5354 = ~n5352 & ~n5353 ;
  assign n5355 = ~n3093 & ~n5354 ;
  assign n5356 = n2989 & ~n5345 ;
  assign n5357 = ~n2989 & ~n5335 ;
  assign n5358 = ~n5356 & ~n5357 ;
  assign n5359 = n3093 & ~n5358 ;
  assign n5360 = ~n5355 & ~n5359 ;
  assign n5361 = ~n3139 & ~n5360 ;
  assign n5362 = ~n5351 & ~n5361 ;
  assign n5363 = ~n3185 & ~n5362 ;
  assign n5364 = x53 & n3185 ;
  assign n5365 = ~n5363 & ~n5364 ;
  assign n5366 = ~n3287 & ~n5365 ;
  assign n5367 = n3093 & ~n5354 ;
  assign n5368 = ~n3093 & ~n5358 ;
  assign n5369 = ~n5367 & ~n5368 ;
  assign n5370 = ~n3242 & ~n5369 ;
  assign n5371 = n3139 & ~n5360 ;
  assign n5372 = ~n3139 & ~n5350 ;
  assign n5373 = ~n5371 & ~n5372 ;
  assign n5374 = n3242 & ~n5373 ;
  assign n5375 = ~n5370 & ~n5374 ;
  assign n5376 = n3287 & ~n5375 ;
  assign n5377 = ~n5366 & ~n5376 ;
  assign n5378 = ~n3335 & ~n5377 ;
  assign n5379 = n3242 & ~n5369 ;
  assign n5380 = ~n3242 & ~n5373 ;
  assign n5381 = ~n5379 & ~n5380 ;
  assign n5382 = n3335 & ~n5381 ;
  assign n5383 = ~n5378 & ~n5382 ;
  assign n5384 = n3484 & ~n5383 ;
  assign n5385 = n3335 & ~n5377 ;
  assign n5386 = ~n3335 & ~n5381 ;
  assign n5387 = ~n5385 & ~n5386 ;
  assign n5388 = n3439 & ~n5387 ;
  assign n5389 = ~n3287 & ~n5375 ;
  assign n5390 = n3287 & ~n5365 ;
  assign n5391 = ~n5389 & ~n5390 ;
  assign n5392 = ~n3384 & ~n5391 ;
  assign n5393 = x21 & n3384 ;
  assign n5394 = ~n5392 & ~n5393 ;
  assign n5395 = ~n3439 & ~n5394 ;
  assign n5396 = ~n5388 & ~n5395 ;
  assign n5397 = ~n3484 & ~n5396 ;
  assign n5398 = ~n5384 & ~n5397 ;
  assign n5399 = x246 & ~n2640 ;
  assign n5400 = x214 & n2640 ;
  assign n5401 = ~n5399 & ~n5400 ;
  assign n5402 = n2693 & ~n5401 ;
  assign n5403 = x182 & ~n2693 ;
  assign n5404 = ~n5402 & ~n5403 ;
  assign n5405 = n2742 & ~n5404 ;
  assign n5406 = x214 & ~n2640 ;
  assign n5407 = x246 & n2640 ;
  assign n5408 = ~n5406 & ~n5407 ;
  assign n5409 = ~n2742 & ~n5408 ;
  assign n5410 = ~n5405 & ~n5409 ;
  assign n5411 = ~n2841 & ~n5410 ;
  assign n5412 = ~n2693 & ~n5401 ;
  assign n5413 = x182 & n2693 ;
  assign n5414 = ~n5412 & ~n5413 ;
  assign n5415 = ~n2791 & ~n5414 ;
  assign n5416 = x150 & n2791 ;
  assign n5417 = ~n5415 & ~n5416 ;
  assign n5418 = n2841 & ~n5417 ;
  assign n5419 = ~n5411 & ~n5418 ;
  assign n5420 = ~n2887 & ~n5419 ;
  assign n5421 = x118 & n2887 ;
  assign n5422 = ~n5420 & ~n5421 ;
  assign n5423 = n2989 & ~n5422 ;
  assign n5424 = n2841 & ~n5410 ;
  assign n5425 = ~n2841 & ~n5417 ;
  assign n5426 = ~n5424 & ~n5425 ;
  assign n5427 = n2944 & ~n5426 ;
  assign n5428 = n2742 & ~n5408 ;
  assign n5429 = ~n2742 & ~n5404 ;
  assign n5430 = ~n5428 & ~n5429 ;
  assign n5431 = ~n2944 & ~n5430 ;
  assign n5432 = ~n5427 & ~n5431 ;
  assign n5433 = ~n2989 & ~n5432 ;
  assign n5434 = ~n5423 & ~n5433 ;
  assign n5435 = ~n3035 & ~n5434 ;
  assign n5436 = x86 & n3035 ;
  assign n5437 = ~n5435 & ~n5436 ;
  assign n5438 = n3139 & ~n5437 ;
  assign n5439 = n2944 & ~n5430 ;
  assign n5440 = ~n2944 & ~n5426 ;
  assign n5441 = ~n5439 & ~n5440 ;
  assign n5442 = ~n3093 & ~n5441 ;
  assign n5443 = n2989 & ~n5432 ;
  assign n5444 = ~n2989 & ~n5422 ;
  assign n5445 = ~n5443 & ~n5444 ;
  assign n5446 = n3093 & ~n5445 ;
  assign n5447 = ~n5442 & ~n5446 ;
  assign n5448 = ~n3139 & ~n5447 ;
  assign n5449 = ~n5438 & ~n5448 ;
  assign n5450 = ~n3185 & ~n5449 ;
  assign n5451 = x54 & n3185 ;
  assign n5452 = ~n5450 & ~n5451 ;
  assign n5453 = ~n3287 & ~n5452 ;
  assign n5454 = n3093 & ~n5441 ;
  assign n5455 = ~n3093 & ~n5445 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = ~n3242 & ~n5456 ;
  assign n5458 = n3139 & ~n5447 ;
  assign n5459 = ~n3139 & ~n5437 ;
  assign n5460 = ~n5458 & ~n5459 ;
  assign n5461 = n3242 & ~n5460 ;
  assign n5462 = ~n5457 & ~n5461 ;
  assign n5463 = n3287 & ~n5462 ;
  assign n5464 = ~n5453 & ~n5463 ;
  assign n5465 = ~n3335 & ~n5464 ;
  assign n5466 = n3242 & ~n5456 ;
  assign n5467 = ~n3242 & ~n5460 ;
  assign n5468 = ~n5466 & ~n5467 ;
  assign n5469 = n3335 & ~n5468 ;
  assign n5470 = ~n5465 & ~n5469 ;
  assign n5471 = n3484 & ~n5470 ;
  assign n5472 = n3335 & ~n5464 ;
  assign n5473 = ~n3335 & ~n5468 ;
  assign n5474 = ~n5472 & ~n5473 ;
  assign n5475 = n3439 & ~n5474 ;
  assign n5476 = ~n3287 & ~n5462 ;
  assign n5477 = n3287 & ~n5452 ;
  assign n5478 = ~n5476 & ~n5477 ;
  assign n5479 = ~n3384 & ~n5478 ;
  assign n5480 = x22 & n3384 ;
  assign n5481 = ~n5479 & ~n5480 ;
  assign n5482 = ~n3439 & ~n5481 ;
  assign n5483 = ~n5475 & ~n5482 ;
  assign n5484 = ~n3484 & ~n5483 ;
  assign n5485 = ~n5471 & ~n5484 ;
  assign n5486 = x247 & ~n2640 ;
  assign n5487 = x215 & n2640 ;
  assign n5488 = ~n5486 & ~n5487 ;
  assign n5489 = n2693 & ~n5488 ;
  assign n5490 = x183 & ~n2693 ;
  assign n5491 = ~n5489 & ~n5490 ;
  assign n5492 = n2742 & ~n5491 ;
  assign n5493 = x215 & ~n2640 ;
  assign n5494 = x247 & n2640 ;
  assign n5495 = ~n5493 & ~n5494 ;
  assign n5496 = ~n2742 & ~n5495 ;
  assign n5497 = ~n5492 & ~n5496 ;
  assign n5498 = ~n2841 & ~n5497 ;
  assign n5499 = ~n2693 & ~n5488 ;
  assign n5500 = x183 & n2693 ;
  assign n5501 = ~n5499 & ~n5500 ;
  assign n5502 = ~n2791 & ~n5501 ;
  assign n5503 = x151 & n2791 ;
  assign n5504 = ~n5502 & ~n5503 ;
  assign n5505 = n2841 & ~n5504 ;
  assign n5506 = ~n5498 & ~n5505 ;
  assign n5507 = ~n2887 & ~n5506 ;
  assign n5508 = x119 & n2887 ;
  assign n5509 = ~n5507 & ~n5508 ;
  assign n5510 = n2989 & ~n5509 ;
  assign n5511 = n2841 & ~n5497 ;
  assign n5512 = ~n2841 & ~n5504 ;
  assign n5513 = ~n5511 & ~n5512 ;
  assign n5514 = n2944 & ~n5513 ;
  assign n5515 = n2742 & ~n5495 ;
  assign n5516 = ~n2742 & ~n5491 ;
  assign n5517 = ~n5515 & ~n5516 ;
  assign n5518 = ~n2944 & ~n5517 ;
  assign n5519 = ~n5514 & ~n5518 ;
  assign n5520 = ~n2989 & ~n5519 ;
  assign n5521 = ~n5510 & ~n5520 ;
  assign n5522 = ~n3035 & ~n5521 ;
  assign n5523 = x87 & n3035 ;
  assign n5524 = ~n5522 & ~n5523 ;
  assign n5525 = n3139 & ~n5524 ;
  assign n5526 = n2944 & ~n5517 ;
  assign n5527 = ~n2944 & ~n5513 ;
  assign n5528 = ~n5526 & ~n5527 ;
  assign n5529 = ~n3093 & ~n5528 ;
  assign n5530 = n2989 & ~n5519 ;
  assign n5531 = ~n2989 & ~n5509 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5533 = n3093 & ~n5532 ;
  assign n5534 = ~n5529 & ~n5533 ;
  assign n5535 = ~n3139 & ~n5534 ;
  assign n5536 = ~n5525 & ~n5535 ;
  assign n5537 = ~n3185 & ~n5536 ;
  assign n5538 = x55 & n3185 ;
  assign n5539 = ~n5537 & ~n5538 ;
  assign n5540 = ~n3287 & ~n5539 ;
  assign n5541 = n3093 & ~n5528 ;
  assign n5542 = ~n3093 & ~n5532 ;
  assign n5543 = ~n5541 & ~n5542 ;
  assign n5544 = ~n3242 & ~n5543 ;
  assign n5545 = n3139 & ~n5534 ;
  assign n5546 = ~n3139 & ~n5524 ;
  assign n5547 = ~n5545 & ~n5546 ;
  assign n5548 = n3242 & ~n5547 ;
  assign n5549 = ~n5544 & ~n5548 ;
  assign n5550 = n3287 & ~n5549 ;
  assign n5551 = ~n5540 & ~n5550 ;
  assign n5552 = ~n3335 & ~n5551 ;
  assign n5553 = n3242 & ~n5543 ;
  assign n5554 = ~n3242 & ~n5547 ;
  assign n5555 = ~n5553 & ~n5554 ;
  assign n5556 = n3335 & ~n5555 ;
  assign n5557 = ~n5552 & ~n5556 ;
  assign n5558 = n3484 & ~n5557 ;
  assign n5559 = n3335 & ~n5551 ;
  assign n5560 = ~n3335 & ~n5555 ;
  assign n5561 = ~n5559 & ~n5560 ;
  assign n5562 = n3439 & ~n5561 ;
  assign n5563 = ~n3287 & ~n5549 ;
  assign n5564 = n3287 & ~n5539 ;
  assign n5565 = ~n5563 & ~n5564 ;
  assign n5566 = ~n3384 & ~n5565 ;
  assign n5567 = x23 & n3384 ;
  assign n5568 = ~n5566 & ~n5567 ;
  assign n5569 = ~n3439 & ~n5568 ;
  assign n5570 = ~n5562 & ~n5569 ;
  assign n5571 = ~n3484 & ~n5570 ;
  assign n5572 = ~n5558 & ~n5571 ;
  assign n5573 = x248 & ~n2640 ;
  assign n5574 = x216 & n2640 ;
  assign n5575 = ~n5573 & ~n5574 ;
  assign n5576 = n2693 & ~n5575 ;
  assign n5577 = x184 & ~n2693 ;
  assign n5578 = ~n5576 & ~n5577 ;
  assign n5579 = n2742 & ~n5578 ;
  assign n5580 = x216 & ~n2640 ;
  assign n5581 = x248 & n2640 ;
  assign n5582 = ~n5580 & ~n5581 ;
  assign n5583 = ~n2742 & ~n5582 ;
  assign n5584 = ~n5579 & ~n5583 ;
  assign n5585 = ~n2841 & ~n5584 ;
  assign n5586 = ~n2693 & ~n5575 ;
  assign n5587 = x184 & n2693 ;
  assign n5588 = ~n5586 & ~n5587 ;
  assign n5589 = ~n2791 & ~n5588 ;
  assign n5590 = x152 & n2791 ;
  assign n5591 = ~n5589 & ~n5590 ;
  assign n5592 = n2841 & ~n5591 ;
  assign n5593 = ~n5585 & ~n5592 ;
  assign n5594 = ~n2887 & ~n5593 ;
  assign n5595 = x120 & n2887 ;
  assign n5596 = ~n5594 & ~n5595 ;
  assign n5597 = n2989 & ~n5596 ;
  assign n5598 = n2841 & ~n5584 ;
  assign n5599 = ~n2841 & ~n5591 ;
  assign n5600 = ~n5598 & ~n5599 ;
  assign n5601 = n2944 & ~n5600 ;
  assign n5602 = n2742 & ~n5582 ;
  assign n5603 = ~n2742 & ~n5578 ;
  assign n5604 = ~n5602 & ~n5603 ;
  assign n5605 = ~n2944 & ~n5604 ;
  assign n5606 = ~n5601 & ~n5605 ;
  assign n5607 = ~n2989 & ~n5606 ;
  assign n5608 = ~n5597 & ~n5607 ;
  assign n5609 = ~n3035 & ~n5608 ;
  assign n5610 = x88 & n3035 ;
  assign n5611 = ~n5609 & ~n5610 ;
  assign n5612 = n3139 & ~n5611 ;
  assign n5613 = n2944 & ~n5604 ;
  assign n5614 = ~n2944 & ~n5600 ;
  assign n5615 = ~n5613 & ~n5614 ;
  assign n5616 = ~n3093 & ~n5615 ;
  assign n5617 = n2989 & ~n5606 ;
  assign n5618 = ~n2989 & ~n5596 ;
  assign n5619 = ~n5617 & ~n5618 ;
  assign n5620 = n3093 & ~n5619 ;
  assign n5621 = ~n5616 & ~n5620 ;
  assign n5622 = ~n3139 & ~n5621 ;
  assign n5623 = ~n5612 & ~n5622 ;
  assign n5624 = ~n3185 & ~n5623 ;
  assign n5625 = x56 & n3185 ;
  assign n5626 = ~n5624 & ~n5625 ;
  assign n5627 = ~n3287 & ~n5626 ;
  assign n5628 = n3093 & ~n5615 ;
  assign n5629 = ~n3093 & ~n5619 ;
  assign n5630 = ~n5628 & ~n5629 ;
  assign n5631 = ~n3242 & ~n5630 ;
  assign n5632 = n3139 & ~n5621 ;
  assign n5633 = ~n3139 & ~n5611 ;
  assign n5634 = ~n5632 & ~n5633 ;
  assign n5635 = n3242 & ~n5634 ;
  assign n5636 = ~n5631 & ~n5635 ;
  assign n5637 = n3287 & ~n5636 ;
  assign n5638 = ~n5627 & ~n5637 ;
  assign n5639 = ~n3335 & ~n5638 ;
  assign n5640 = n3242 & ~n5630 ;
  assign n5641 = ~n3242 & ~n5634 ;
  assign n5642 = ~n5640 & ~n5641 ;
  assign n5643 = n3335 & ~n5642 ;
  assign n5644 = ~n5639 & ~n5643 ;
  assign n5645 = n3484 & ~n5644 ;
  assign n5646 = n3335 & ~n5638 ;
  assign n5647 = ~n3335 & ~n5642 ;
  assign n5648 = ~n5646 & ~n5647 ;
  assign n5649 = n3439 & ~n5648 ;
  assign n5650 = ~n3287 & ~n5636 ;
  assign n5651 = n3287 & ~n5626 ;
  assign n5652 = ~n5650 & ~n5651 ;
  assign n5653 = ~n3384 & ~n5652 ;
  assign n5654 = x24 & n3384 ;
  assign n5655 = ~n5653 & ~n5654 ;
  assign n5656 = ~n3439 & ~n5655 ;
  assign n5657 = ~n5649 & ~n5656 ;
  assign n5658 = ~n3484 & ~n5657 ;
  assign n5659 = ~n5645 & ~n5658 ;
  assign n5660 = x249 & ~n2640 ;
  assign n5661 = x217 & n2640 ;
  assign n5662 = ~n5660 & ~n5661 ;
  assign n5663 = n2693 & ~n5662 ;
  assign n5664 = x185 & ~n2693 ;
  assign n5665 = ~n5663 & ~n5664 ;
  assign n5666 = n2742 & ~n5665 ;
  assign n5667 = x217 & ~n2640 ;
  assign n5668 = x249 & n2640 ;
  assign n5669 = ~n5667 & ~n5668 ;
  assign n5670 = ~n2742 & ~n5669 ;
  assign n5671 = ~n5666 & ~n5670 ;
  assign n5672 = ~n2841 & ~n5671 ;
  assign n5673 = ~n2693 & ~n5662 ;
  assign n5674 = x185 & n2693 ;
  assign n5675 = ~n5673 & ~n5674 ;
  assign n5676 = ~n2791 & ~n5675 ;
  assign n5677 = x153 & n2791 ;
  assign n5678 = ~n5676 & ~n5677 ;
  assign n5679 = n2841 & ~n5678 ;
  assign n5680 = ~n5672 & ~n5679 ;
  assign n5681 = ~n2887 & ~n5680 ;
  assign n5682 = x121 & n2887 ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5684 = n2989 & ~n5683 ;
  assign n5685 = n2841 & ~n5671 ;
  assign n5686 = ~n2841 & ~n5678 ;
  assign n5687 = ~n5685 & ~n5686 ;
  assign n5688 = n2944 & ~n5687 ;
  assign n5689 = n2742 & ~n5669 ;
  assign n5690 = ~n2742 & ~n5665 ;
  assign n5691 = ~n5689 & ~n5690 ;
  assign n5692 = ~n2944 & ~n5691 ;
  assign n5693 = ~n5688 & ~n5692 ;
  assign n5694 = ~n2989 & ~n5693 ;
  assign n5695 = ~n5684 & ~n5694 ;
  assign n5696 = ~n3035 & ~n5695 ;
  assign n5697 = x89 & n3035 ;
  assign n5698 = ~n5696 & ~n5697 ;
  assign n5699 = n3139 & ~n5698 ;
  assign n5700 = n2944 & ~n5691 ;
  assign n5701 = ~n2944 & ~n5687 ;
  assign n5702 = ~n5700 & ~n5701 ;
  assign n5703 = ~n3093 & ~n5702 ;
  assign n5704 = n2989 & ~n5693 ;
  assign n5705 = ~n2989 & ~n5683 ;
  assign n5706 = ~n5704 & ~n5705 ;
  assign n5707 = n3093 & ~n5706 ;
  assign n5708 = ~n5703 & ~n5707 ;
  assign n5709 = ~n3139 & ~n5708 ;
  assign n5710 = ~n5699 & ~n5709 ;
  assign n5711 = ~n3185 & ~n5710 ;
  assign n5712 = x57 & n3185 ;
  assign n5713 = ~n5711 & ~n5712 ;
  assign n5714 = ~n3287 & ~n5713 ;
  assign n5715 = n3093 & ~n5702 ;
  assign n5716 = ~n3093 & ~n5706 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = ~n3242 & ~n5717 ;
  assign n5719 = n3139 & ~n5708 ;
  assign n5720 = ~n3139 & ~n5698 ;
  assign n5721 = ~n5719 & ~n5720 ;
  assign n5722 = n3242 & ~n5721 ;
  assign n5723 = ~n5718 & ~n5722 ;
  assign n5724 = n3287 & ~n5723 ;
  assign n5725 = ~n5714 & ~n5724 ;
  assign n5726 = ~n3335 & ~n5725 ;
  assign n5727 = n3242 & ~n5717 ;
  assign n5728 = ~n3242 & ~n5721 ;
  assign n5729 = ~n5727 & ~n5728 ;
  assign n5730 = n3335 & ~n5729 ;
  assign n5731 = ~n5726 & ~n5730 ;
  assign n5732 = n3484 & ~n5731 ;
  assign n5733 = n3335 & ~n5725 ;
  assign n5734 = ~n3335 & ~n5729 ;
  assign n5735 = ~n5733 & ~n5734 ;
  assign n5736 = n3439 & ~n5735 ;
  assign n5737 = ~n3287 & ~n5723 ;
  assign n5738 = n3287 & ~n5713 ;
  assign n5739 = ~n5737 & ~n5738 ;
  assign n5740 = ~n3384 & ~n5739 ;
  assign n5741 = x25 & n3384 ;
  assign n5742 = ~n5740 & ~n5741 ;
  assign n5743 = ~n3439 & ~n5742 ;
  assign n5744 = ~n5736 & ~n5743 ;
  assign n5745 = ~n3484 & ~n5744 ;
  assign n5746 = ~n5732 & ~n5745 ;
  assign n5747 = x250 & ~n2640 ;
  assign n5748 = x218 & n2640 ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5750 = n2693 & ~n5749 ;
  assign n5751 = x186 & ~n2693 ;
  assign n5752 = ~n5750 & ~n5751 ;
  assign n5753 = n2742 & ~n5752 ;
  assign n5754 = x218 & ~n2640 ;
  assign n5755 = x250 & n2640 ;
  assign n5756 = ~n5754 & ~n5755 ;
  assign n5757 = ~n2742 & ~n5756 ;
  assign n5758 = ~n5753 & ~n5757 ;
  assign n5759 = ~n2841 & ~n5758 ;
  assign n5760 = ~n2693 & ~n5749 ;
  assign n5761 = x186 & n2693 ;
  assign n5762 = ~n5760 & ~n5761 ;
  assign n5763 = ~n2791 & ~n5762 ;
  assign n5764 = x154 & n2791 ;
  assign n5765 = ~n5763 & ~n5764 ;
  assign n5766 = n2841 & ~n5765 ;
  assign n5767 = ~n5759 & ~n5766 ;
  assign n5768 = ~n2887 & ~n5767 ;
  assign n5769 = x122 & n2887 ;
  assign n5770 = ~n5768 & ~n5769 ;
  assign n5771 = n2989 & ~n5770 ;
  assign n5772 = n2841 & ~n5758 ;
  assign n5773 = ~n2841 & ~n5765 ;
  assign n5774 = ~n5772 & ~n5773 ;
  assign n5775 = n2944 & ~n5774 ;
  assign n5776 = n2742 & ~n5756 ;
  assign n5777 = ~n2742 & ~n5752 ;
  assign n5778 = ~n5776 & ~n5777 ;
  assign n5779 = ~n2944 & ~n5778 ;
  assign n5780 = ~n5775 & ~n5779 ;
  assign n5781 = ~n2989 & ~n5780 ;
  assign n5782 = ~n5771 & ~n5781 ;
  assign n5783 = ~n3035 & ~n5782 ;
  assign n5784 = x90 & n3035 ;
  assign n5785 = ~n5783 & ~n5784 ;
  assign n5786 = n3139 & ~n5785 ;
  assign n5787 = n2944 & ~n5778 ;
  assign n5788 = ~n2944 & ~n5774 ;
  assign n5789 = ~n5787 & ~n5788 ;
  assign n5790 = ~n3093 & ~n5789 ;
  assign n5791 = n2989 & ~n5780 ;
  assign n5792 = ~n2989 & ~n5770 ;
  assign n5793 = ~n5791 & ~n5792 ;
  assign n5794 = n3093 & ~n5793 ;
  assign n5795 = ~n5790 & ~n5794 ;
  assign n5796 = ~n3139 & ~n5795 ;
  assign n5797 = ~n5786 & ~n5796 ;
  assign n5798 = ~n3185 & ~n5797 ;
  assign n5799 = x58 & n3185 ;
  assign n5800 = ~n5798 & ~n5799 ;
  assign n5801 = ~n3287 & ~n5800 ;
  assign n5802 = n3093 & ~n5789 ;
  assign n5803 = ~n3093 & ~n5793 ;
  assign n5804 = ~n5802 & ~n5803 ;
  assign n5805 = ~n3242 & ~n5804 ;
  assign n5806 = n3139 & ~n5795 ;
  assign n5807 = ~n3139 & ~n5785 ;
  assign n5808 = ~n5806 & ~n5807 ;
  assign n5809 = n3242 & ~n5808 ;
  assign n5810 = ~n5805 & ~n5809 ;
  assign n5811 = n3287 & ~n5810 ;
  assign n5812 = ~n5801 & ~n5811 ;
  assign n5813 = ~n3335 & ~n5812 ;
  assign n5814 = n3242 & ~n5804 ;
  assign n5815 = ~n3242 & ~n5808 ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = n3335 & ~n5816 ;
  assign n5818 = ~n5813 & ~n5817 ;
  assign n5819 = n3484 & ~n5818 ;
  assign n5820 = n3335 & ~n5812 ;
  assign n5821 = ~n3335 & ~n5816 ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5823 = n3439 & ~n5822 ;
  assign n5824 = ~n3287 & ~n5810 ;
  assign n5825 = n3287 & ~n5800 ;
  assign n5826 = ~n5824 & ~n5825 ;
  assign n5827 = ~n3384 & ~n5826 ;
  assign n5828 = x26 & n3384 ;
  assign n5829 = ~n5827 & ~n5828 ;
  assign n5830 = ~n3439 & ~n5829 ;
  assign n5831 = ~n5823 & ~n5830 ;
  assign n5832 = ~n3484 & ~n5831 ;
  assign n5833 = ~n5819 & ~n5832 ;
  assign n5834 = x251 & ~n2640 ;
  assign n5835 = x219 & n2640 ;
  assign n5836 = ~n5834 & ~n5835 ;
  assign n5837 = n2693 & ~n5836 ;
  assign n5838 = x187 & ~n2693 ;
  assign n5839 = ~n5837 & ~n5838 ;
  assign n5840 = n2742 & ~n5839 ;
  assign n5841 = x219 & ~n2640 ;
  assign n5842 = x251 & n2640 ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = ~n2742 & ~n5843 ;
  assign n5845 = ~n5840 & ~n5844 ;
  assign n5846 = ~n2841 & ~n5845 ;
  assign n5847 = ~n2693 & ~n5836 ;
  assign n5848 = x187 & n2693 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = ~n2791 & ~n5849 ;
  assign n5851 = x155 & n2791 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = n2841 & ~n5852 ;
  assign n5854 = ~n5846 & ~n5853 ;
  assign n5855 = ~n2887 & ~n5854 ;
  assign n5856 = x123 & n2887 ;
  assign n5857 = ~n5855 & ~n5856 ;
  assign n5858 = n2989 & ~n5857 ;
  assign n5859 = n2841 & ~n5845 ;
  assign n5860 = ~n2841 & ~n5852 ;
  assign n5861 = ~n5859 & ~n5860 ;
  assign n5862 = n2944 & ~n5861 ;
  assign n5863 = n2742 & ~n5843 ;
  assign n5864 = ~n2742 & ~n5839 ;
  assign n5865 = ~n5863 & ~n5864 ;
  assign n5866 = ~n2944 & ~n5865 ;
  assign n5867 = ~n5862 & ~n5866 ;
  assign n5868 = ~n2989 & ~n5867 ;
  assign n5869 = ~n5858 & ~n5868 ;
  assign n5870 = ~n3035 & ~n5869 ;
  assign n5871 = x91 & n3035 ;
  assign n5872 = ~n5870 & ~n5871 ;
  assign n5873 = n3139 & ~n5872 ;
  assign n5874 = n2944 & ~n5865 ;
  assign n5875 = ~n2944 & ~n5861 ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = ~n3093 & ~n5876 ;
  assign n5878 = n2989 & ~n5867 ;
  assign n5879 = ~n2989 & ~n5857 ;
  assign n5880 = ~n5878 & ~n5879 ;
  assign n5881 = n3093 & ~n5880 ;
  assign n5882 = ~n5877 & ~n5881 ;
  assign n5883 = ~n3139 & ~n5882 ;
  assign n5884 = ~n5873 & ~n5883 ;
  assign n5885 = ~n3185 & ~n5884 ;
  assign n5886 = x59 & n3185 ;
  assign n5887 = ~n5885 & ~n5886 ;
  assign n5888 = ~n3287 & ~n5887 ;
  assign n5889 = n3093 & ~n5876 ;
  assign n5890 = ~n3093 & ~n5880 ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = ~n3242 & ~n5891 ;
  assign n5893 = n3139 & ~n5882 ;
  assign n5894 = ~n3139 & ~n5872 ;
  assign n5895 = ~n5893 & ~n5894 ;
  assign n5896 = n3242 & ~n5895 ;
  assign n5897 = ~n5892 & ~n5896 ;
  assign n5898 = n3287 & ~n5897 ;
  assign n5899 = ~n5888 & ~n5898 ;
  assign n5900 = ~n3335 & ~n5899 ;
  assign n5901 = n3242 & ~n5891 ;
  assign n5902 = ~n3242 & ~n5895 ;
  assign n5903 = ~n5901 & ~n5902 ;
  assign n5904 = n3335 & ~n5903 ;
  assign n5905 = ~n5900 & ~n5904 ;
  assign n5906 = n3484 & ~n5905 ;
  assign n5907 = n3335 & ~n5899 ;
  assign n5908 = ~n3335 & ~n5903 ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = n3439 & ~n5909 ;
  assign n5911 = ~n3287 & ~n5897 ;
  assign n5912 = n3287 & ~n5887 ;
  assign n5913 = ~n5911 & ~n5912 ;
  assign n5914 = ~n3384 & ~n5913 ;
  assign n5915 = x27 & n3384 ;
  assign n5916 = ~n5914 & ~n5915 ;
  assign n5917 = ~n3439 & ~n5916 ;
  assign n5918 = ~n5910 & ~n5917 ;
  assign n5919 = ~n3484 & ~n5918 ;
  assign n5920 = ~n5906 & ~n5919 ;
  assign n5921 = x252 & ~n2640 ;
  assign n5922 = x220 & n2640 ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5924 = n2693 & ~n5923 ;
  assign n5925 = x188 & ~n2693 ;
  assign n5926 = ~n5924 & ~n5925 ;
  assign n5927 = n2742 & ~n5926 ;
  assign n5928 = x220 & ~n2640 ;
  assign n5929 = x252 & n2640 ;
  assign n5930 = ~n5928 & ~n5929 ;
  assign n5931 = ~n2742 & ~n5930 ;
  assign n5932 = ~n5927 & ~n5931 ;
  assign n5933 = ~n2841 & ~n5932 ;
  assign n5934 = ~n2693 & ~n5923 ;
  assign n5935 = x188 & n2693 ;
  assign n5936 = ~n5934 & ~n5935 ;
  assign n5937 = ~n2791 & ~n5936 ;
  assign n5938 = x156 & n2791 ;
  assign n5939 = ~n5937 & ~n5938 ;
  assign n5940 = n2841 & ~n5939 ;
  assign n5941 = ~n5933 & ~n5940 ;
  assign n5942 = ~n2887 & ~n5941 ;
  assign n5943 = x124 & n2887 ;
  assign n5944 = ~n5942 & ~n5943 ;
  assign n5945 = n2989 & ~n5944 ;
  assign n5946 = n2841 & ~n5932 ;
  assign n5947 = ~n2841 & ~n5939 ;
  assign n5948 = ~n5946 & ~n5947 ;
  assign n5949 = n2944 & ~n5948 ;
  assign n5950 = n2742 & ~n5930 ;
  assign n5951 = ~n2742 & ~n5926 ;
  assign n5952 = ~n5950 & ~n5951 ;
  assign n5953 = ~n2944 & ~n5952 ;
  assign n5954 = ~n5949 & ~n5953 ;
  assign n5955 = ~n2989 & ~n5954 ;
  assign n5956 = ~n5945 & ~n5955 ;
  assign n5957 = ~n3035 & ~n5956 ;
  assign n5958 = x92 & n3035 ;
  assign n5959 = ~n5957 & ~n5958 ;
  assign n5960 = n3139 & ~n5959 ;
  assign n5961 = n2944 & ~n5952 ;
  assign n5962 = ~n2944 & ~n5948 ;
  assign n5963 = ~n5961 & ~n5962 ;
  assign n5964 = ~n3093 & ~n5963 ;
  assign n5965 = n2989 & ~n5954 ;
  assign n5966 = ~n2989 & ~n5944 ;
  assign n5967 = ~n5965 & ~n5966 ;
  assign n5968 = n3093 & ~n5967 ;
  assign n5969 = ~n5964 & ~n5968 ;
  assign n5970 = ~n3139 & ~n5969 ;
  assign n5971 = ~n5960 & ~n5970 ;
  assign n5972 = ~n3185 & ~n5971 ;
  assign n5973 = x60 & n3185 ;
  assign n5974 = ~n5972 & ~n5973 ;
  assign n5975 = ~n3287 & ~n5974 ;
  assign n5976 = n3093 & ~n5963 ;
  assign n5977 = ~n3093 & ~n5967 ;
  assign n5978 = ~n5976 & ~n5977 ;
  assign n5979 = ~n3242 & ~n5978 ;
  assign n5980 = n3139 & ~n5969 ;
  assign n5981 = ~n3139 & ~n5959 ;
  assign n5982 = ~n5980 & ~n5981 ;
  assign n5983 = n3242 & ~n5982 ;
  assign n5984 = ~n5979 & ~n5983 ;
  assign n5985 = n3287 & ~n5984 ;
  assign n5986 = ~n5975 & ~n5985 ;
  assign n5987 = ~n3335 & ~n5986 ;
  assign n5988 = n3242 & ~n5978 ;
  assign n5989 = ~n3242 & ~n5982 ;
  assign n5990 = ~n5988 & ~n5989 ;
  assign n5991 = n3335 & ~n5990 ;
  assign n5992 = ~n5987 & ~n5991 ;
  assign n5993 = n3484 & ~n5992 ;
  assign n5994 = n3335 & ~n5986 ;
  assign n5995 = ~n3335 & ~n5990 ;
  assign n5996 = ~n5994 & ~n5995 ;
  assign n5997 = n3439 & ~n5996 ;
  assign n5998 = ~n3287 & ~n5984 ;
  assign n5999 = n3287 & ~n5974 ;
  assign n6000 = ~n5998 & ~n5999 ;
  assign n6001 = ~n3384 & ~n6000 ;
  assign n6002 = x28 & n3384 ;
  assign n6003 = ~n6001 & ~n6002 ;
  assign n6004 = ~n3439 & ~n6003 ;
  assign n6005 = ~n5997 & ~n6004 ;
  assign n6006 = ~n3484 & ~n6005 ;
  assign n6007 = ~n5993 & ~n6006 ;
  assign n6008 = x253 & ~n2640 ;
  assign n6009 = x221 & n2640 ;
  assign n6010 = ~n6008 & ~n6009 ;
  assign n6011 = n2693 & ~n6010 ;
  assign n6012 = x189 & ~n2693 ;
  assign n6013 = ~n6011 & ~n6012 ;
  assign n6014 = n2742 & ~n6013 ;
  assign n6015 = x221 & ~n2640 ;
  assign n6016 = x253 & n2640 ;
  assign n6017 = ~n6015 & ~n6016 ;
  assign n6018 = ~n2742 & ~n6017 ;
  assign n6019 = ~n6014 & ~n6018 ;
  assign n6020 = ~n2841 & ~n6019 ;
  assign n6021 = ~n2693 & ~n6010 ;
  assign n6022 = x189 & n2693 ;
  assign n6023 = ~n6021 & ~n6022 ;
  assign n6024 = ~n2791 & ~n6023 ;
  assign n6025 = x157 & n2791 ;
  assign n6026 = ~n6024 & ~n6025 ;
  assign n6027 = n2841 & ~n6026 ;
  assign n6028 = ~n6020 & ~n6027 ;
  assign n6029 = ~n2887 & ~n6028 ;
  assign n6030 = x125 & n2887 ;
  assign n6031 = ~n6029 & ~n6030 ;
  assign n6032 = n2989 & ~n6031 ;
  assign n6033 = n2841 & ~n6019 ;
  assign n6034 = ~n2841 & ~n6026 ;
  assign n6035 = ~n6033 & ~n6034 ;
  assign n6036 = n2944 & ~n6035 ;
  assign n6037 = n2742 & ~n6017 ;
  assign n6038 = ~n2742 & ~n6013 ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6040 = ~n2944 & ~n6039 ;
  assign n6041 = ~n6036 & ~n6040 ;
  assign n6042 = ~n2989 & ~n6041 ;
  assign n6043 = ~n6032 & ~n6042 ;
  assign n6044 = ~n3035 & ~n6043 ;
  assign n6045 = x93 & n3035 ;
  assign n6046 = ~n6044 & ~n6045 ;
  assign n6047 = n3139 & ~n6046 ;
  assign n6048 = n2944 & ~n6039 ;
  assign n6049 = ~n2944 & ~n6035 ;
  assign n6050 = ~n6048 & ~n6049 ;
  assign n6051 = ~n3093 & ~n6050 ;
  assign n6052 = n2989 & ~n6041 ;
  assign n6053 = ~n2989 & ~n6031 ;
  assign n6054 = ~n6052 & ~n6053 ;
  assign n6055 = n3093 & ~n6054 ;
  assign n6056 = ~n6051 & ~n6055 ;
  assign n6057 = ~n3139 & ~n6056 ;
  assign n6058 = ~n6047 & ~n6057 ;
  assign n6059 = ~n3185 & ~n6058 ;
  assign n6060 = x61 & n3185 ;
  assign n6061 = ~n6059 & ~n6060 ;
  assign n6062 = ~n3287 & ~n6061 ;
  assign n6063 = n3093 & ~n6050 ;
  assign n6064 = ~n3093 & ~n6054 ;
  assign n6065 = ~n6063 & ~n6064 ;
  assign n6066 = ~n3242 & ~n6065 ;
  assign n6067 = n3139 & ~n6056 ;
  assign n6068 = ~n3139 & ~n6046 ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6070 = n3242 & ~n6069 ;
  assign n6071 = ~n6066 & ~n6070 ;
  assign n6072 = n3287 & ~n6071 ;
  assign n6073 = ~n6062 & ~n6072 ;
  assign n6074 = ~n3335 & ~n6073 ;
  assign n6075 = n3242 & ~n6065 ;
  assign n6076 = ~n3242 & ~n6069 ;
  assign n6077 = ~n6075 & ~n6076 ;
  assign n6078 = n3335 & ~n6077 ;
  assign n6079 = ~n6074 & ~n6078 ;
  assign n6080 = n3484 & ~n6079 ;
  assign n6081 = n3335 & ~n6073 ;
  assign n6082 = ~n3335 & ~n6077 ;
  assign n6083 = ~n6081 & ~n6082 ;
  assign n6084 = n3439 & ~n6083 ;
  assign n6085 = ~n3287 & ~n6071 ;
  assign n6086 = n3287 & ~n6061 ;
  assign n6087 = ~n6085 & ~n6086 ;
  assign n6088 = ~n3384 & ~n6087 ;
  assign n6089 = x29 & n3384 ;
  assign n6090 = ~n6088 & ~n6089 ;
  assign n6091 = ~n3439 & ~n6090 ;
  assign n6092 = ~n6084 & ~n6091 ;
  assign n6093 = ~n3484 & ~n6092 ;
  assign n6094 = ~n6080 & ~n6093 ;
  assign n6095 = x254 & ~n2640 ;
  assign n6096 = x222 & n2640 ;
  assign n6097 = ~n6095 & ~n6096 ;
  assign n6098 = n2693 & ~n6097 ;
  assign n6099 = x190 & ~n2693 ;
  assign n6100 = ~n6098 & ~n6099 ;
  assign n6101 = n2742 & ~n6100 ;
  assign n6102 = x222 & ~n2640 ;
  assign n6103 = x254 & n2640 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6105 = ~n2742 & ~n6104 ;
  assign n6106 = ~n6101 & ~n6105 ;
  assign n6107 = ~n2841 & ~n6106 ;
  assign n6108 = ~n2693 & ~n6097 ;
  assign n6109 = x190 & n2693 ;
  assign n6110 = ~n6108 & ~n6109 ;
  assign n6111 = ~n2791 & ~n6110 ;
  assign n6112 = x158 & n2791 ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = n2841 & ~n6113 ;
  assign n6115 = ~n6107 & ~n6114 ;
  assign n6116 = ~n2887 & ~n6115 ;
  assign n6117 = x126 & n2887 ;
  assign n6118 = ~n6116 & ~n6117 ;
  assign n6119 = n2989 & ~n6118 ;
  assign n6120 = n2841 & ~n6106 ;
  assign n6121 = ~n2841 & ~n6113 ;
  assign n6122 = ~n6120 & ~n6121 ;
  assign n6123 = n2944 & ~n6122 ;
  assign n6124 = n2742 & ~n6104 ;
  assign n6125 = ~n2742 & ~n6100 ;
  assign n6126 = ~n6124 & ~n6125 ;
  assign n6127 = ~n2944 & ~n6126 ;
  assign n6128 = ~n6123 & ~n6127 ;
  assign n6129 = ~n2989 & ~n6128 ;
  assign n6130 = ~n6119 & ~n6129 ;
  assign n6131 = ~n3035 & ~n6130 ;
  assign n6132 = x94 & n3035 ;
  assign n6133 = ~n6131 & ~n6132 ;
  assign n6134 = n3139 & ~n6133 ;
  assign n6135 = n2944 & ~n6126 ;
  assign n6136 = ~n2944 & ~n6122 ;
  assign n6137 = ~n6135 & ~n6136 ;
  assign n6138 = ~n3093 & ~n6137 ;
  assign n6139 = n2989 & ~n6128 ;
  assign n6140 = ~n2989 & ~n6118 ;
  assign n6141 = ~n6139 & ~n6140 ;
  assign n6142 = n3093 & ~n6141 ;
  assign n6143 = ~n6138 & ~n6142 ;
  assign n6144 = ~n3139 & ~n6143 ;
  assign n6145 = ~n6134 & ~n6144 ;
  assign n6146 = ~n3185 & ~n6145 ;
  assign n6147 = x62 & n3185 ;
  assign n6148 = ~n6146 & ~n6147 ;
  assign n6149 = ~n3287 & ~n6148 ;
  assign n6150 = n3093 & ~n6137 ;
  assign n6151 = ~n3093 & ~n6141 ;
  assign n6152 = ~n6150 & ~n6151 ;
  assign n6153 = ~n3242 & ~n6152 ;
  assign n6154 = n3139 & ~n6143 ;
  assign n6155 = ~n3139 & ~n6133 ;
  assign n6156 = ~n6154 & ~n6155 ;
  assign n6157 = n3242 & ~n6156 ;
  assign n6158 = ~n6153 & ~n6157 ;
  assign n6159 = n3287 & ~n6158 ;
  assign n6160 = ~n6149 & ~n6159 ;
  assign n6161 = ~n3335 & ~n6160 ;
  assign n6162 = n3242 & ~n6152 ;
  assign n6163 = ~n3242 & ~n6156 ;
  assign n6164 = ~n6162 & ~n6163 ;
  assign n6165 = n3335 & ~n6164 ;
  assign n6166 = ~n6161 & ~n6165 ;
  assign n6167 = n3484 & ~n6166 ;
  assign n6168 = n3335 & ~n6160 ;
  assign n6169 = ~n3335 & ~n6164 ;
  assign n6170 = ~n6168 & ~n6169 ;
  assign n6171 = n3439 & ~n6170 ;
  assign n6172 = ~n3287 & ~n6158 ;
  assign n6173 = n3287 & ~n6148 ;
  assign n6174 = ~n6172 & ~n6173 ;
  assign n6175 = ~n3384 & ~n6174 ;
  assign n6176 = x30 & n3384 ;
  assign n6177 = ~n6175 & ~n6176 ;
  assign n6178 = ~n3439 & ~n6177 ;
  assign n6179 = ~n6171 & ~n6178 ;
  assign n6180 = ~n3484 & ~n6179 ;
  assign n6181 = ~n6167 & ~n6180 ;
  assign n6182 = x255 & ~n2640 ;
  assign n6183 = x223 & n2640 ;
  assign n6184 = ~n6182 & ~n6183 ;
  assign n6185 = n2693 & ~n6184 ;
  assign n6186 = x191 & ~n2693 ;
  assign n6187 = ~n6185 & ~n6186 ;
  assign n6188 = n2742 & ~n6187 ;
  assign n6189 = x223 & ~n2640 ;
  assign n6190 = x255 & n2640 ;
  assign n6191 = ~n6189 & ~n6190 ;
  assign n6192 = ~n2742 & ~n6191 ;
  assign n6193 = ~n6188 & ~n6192 ;
  assign n6194 = ~n2841 & ~n6193 ;
  assign n6195 = ~n2693 & ~n6184 ;
  assign n6196 = x191 & n2693 ;
  assign n6197 = ~n6195 & ~n6196 ;
  assign n6198 = ~n2791 & ~n6197 ;
  assign n6199 = x159 & n2791 ;
  assign n6200 = ~n6198 & ~n6199 ;
  assign n6201 = n2841 & ~n6200 ;
  assign n6202 = ~n6194 & ~n6201 ;
  assign n6203 = ~n2887 & ~n6202 ;
  assign n6204 = x127 & n2887 ;
  assign n6205 = ~n6203 & ~n6204 ;
  assign n6206 = n2989 & ~n6205 ;
  assign n6207 = n2841 & ~n6193 ;
  assign n6208 = ~n2841 & ~n6200 ;
  assign n6209 = ~n6207 & ~n6208 ;
  assign n6210 = n2944 & ~n6209 ;
  assign n6211 = n2742 & ~n6191 ;
  assign n6212 = ~n2742 & ~n6187 ;
  assign n6213 = ~n6211 & ~n6212 ;
  assign n6214 = ~n2944 & ~n6213 ;
  assign n6215 = ~n6210 & ~n6214 ;
  assign n6216 = ~n2989 & ~n6215 ;
  assign n6217 = ~n6206 & ~n6216 ;
  assign n6218 = ~n3035 & ~n6217 ;
  assign n6219 = x95 & n3035 ;
  assign n6220 = ~n6218 & ~n6219 ;
  assign n6221 = n3139 & ~n6220 ;
  assign n6222 = n2944 & ~n6213 ;
  assign n6223 = ~n2944 & ~n6209 ;
  assign n6224 = ~n6222 & ~n6223 ;
  assign n6225 = ~n3093 & ~n6224 ;
  assign n6226 = n2989 & ~n6215 ;
  assign n6227 = ~n2989 & ~n6205 ;
  assign n6228 = ~n6226 & ~n6227 ;
  assign n6229 = n3093 & ~n6228 ;
  assign n6230 = ~n6225 & ~n6229 ;
  assign n6231 = ~n3139 & ~n6230 ;
  assign n6232 = ~n6221 & ~n6231 ;
  assign n6233 = ~n3185 & ~n6232 ;
  assign n6234 = x63 & n3185 ;
  assign n6235 = ~n6233 & ~n6234 ;
  assign n6236 = ~n3287 & ~n6235 ;
  assign n6237 = n3093 & ~n6224 ;
  assign n6238 = ~n3093 & ~n6228 ;
  assign n6239 = ~n6237 & ~n6238 ;
  assign n6240 = ~n3242 & ~n6239 ;
  assign n6241 = n3139 & ~n6230 ;
  assign n6242 = ~n3139 & ~n6220 ;
  assign n6243 = ~n6241 & ~n6242 ;
  assign n6244 = n3242 & ~n6243 ;
  assign n6245 = ~n6240 & ~n6244 ;
  assign n6246 = n3287 & ~n6245 ;
  assign n6247 = ~n6236 & ~n6246 ;
  assign n6248 = ~n3335 & ~n6247 ;
  assign n6249 = n3242 & ~n6239 ;
  assign n6250 = ~n3242 & ~n6243 ;
  assign n6251 = ~n6249 & ~n6250 ;
  assign n6252 = n3335 & ~n6251 ;
  assign n6253 = ~n6248 & ~n6252 ;
  assign n6254 = n3484 & ~n6253 ;
  assign n6255 = n3335 & ~n6247 ;
  assign n6256 = ~n3335 & ~n6251 ;
  assign n6257 = ~n6255 & ~n6256 ;
  assign n6258 = n3439 & ~n6257 ;
  assign n6259 = ~n3287 & ~n6245 ;
  assign n6260 = n3287 & ~n6235 ;
  assign n6261 = ~n6259 & ~n6260 ;
  assign n6262 = ~n3384 & ~n6261 ;
  assign n6263 = x31 & n3384 ;
  assign n6264 = ~n6262 & ~n6263 ;
  assign n6265 = ~n3439 & ~n6264 ;
  assign n6266 = ~n6258 & ~n6265 ;
  assign n6267 = ~n3484 & ~n6266 ;
  assign n6268 = ~n6254 & ~n6267 ;
  assign n6269 = ~n3484 & ~n3569 ;
  assign n6270 = n3484 & ~n3565 ;
  assign n6271 = ~n6269 & ~n6270 ;
  assign n6272 = ~n3484 & ~n3643 ;
  assign n6273 = n3484 & ~n3656 ;
  assign n6274 = ~n6272 & ~n6273 ;
  assign n6275 = ~n3484 & ~n3730 ;
  assign n6276 = n3484 & ~n3743 ;
  assign n6277 = ~n6275 & ~n6276 ;
  assign n6278 = ~n3484 & ~n3817 ;
  assign n6279 = n3484 & ~n3830 ;
  assign n6280 = ~n6278 & ~n6279 ;
  assign n6281 = ~n3484 & ~n3904 ;
  assign n6282 = n3484 & ~n3917 ;
  assign n6283 = ~n6281 & ~n6282 ;
  assign n6284 = ~n3484 & ~n3991 ;
  assign n6285 = n3484 & ~n4004 ;
  assign n6286 = ~n6284 & ~n6285 ;
  assign n6287 = ~n3484 & ~n4078 ;
  assign n6288 = n3484 & ~n4091 ;
  assign n6289 = ~n6287 & ~n6288 ;
  assign n6290 = ~n3484 & ~n4165 ;
  assign n6291 = n3484 & ~n4178 ;
  assign n6292 = ~n6290 & ~n6291 ;
  assign n6293 = ~n3484 & ~n4252 ;
  assign n6294 = n3484 & ~n4265 ;
  assign n6295 = ~n6293 & ~n6294 ;
  assign n6296 = ~n3484 & ~n4339 ;
  assign n6297 = n3484 & ~n4352 ;
  assign n6298 = ~n6296 & ~n6297 ;
  assign n6299 = ~n3484 & ~n4426 ;
  assign n6300 = n3484 & ~n4439 ;
  assign n6301 = ~n6299 & ~n6300 ;
  assign n6302 = ~n3484 & ~n4513 ;
  assign n6303 = n3484 & ~n4526 ;
  assign n6304 = ~n6302 & ~n6303 ;
  assign n6305 = ~n3484 & ~n4600 ;
  assign n6306 = n3484 & ~n4613 ;
  assign n6307 = ~n6305 & ~n6306 ;
  assign n6308 = ~n3484 & ~n4687 ;
  assign n6309 = n3484 & ~n4700 ;
  assign n6310 = ~n6308 & ~n6309 ;
  assign n6311 = ~n3484 & ~n4774 ;
  assign n6312 = n3484 & ~n4787 ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = ~n3484 & ~n4861 ;
  assign n6315 = n3484 & ~n4874 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = ~n3484 & ~n4948 ;
  assign n6318 = n3484 & ~n4961 ;
  assign n6319 = ~n6317 & ~n6318 ;
  assign n6320 = ~n3484 & ~n5035 ;
  assign n6321 = n3484 & ~n5048 ;
  assign n6322 = ~n6320 & ~n6321 ;
  assign n6323 = ~n3484 & ~n5122 ;
  assign n6324 = n3484 & ~n5135 ;
  assign n6325 = ~n6323 & ~n6324 ;
  assign n6326 = ~n3484 & ~n5209 ;
  assign n6327 = n3484 & ~n5222 ;
  assign n6328 = ~n6326 & ~n6327 ;
  assign n6329 = ~n3484 & ~n5296 ;
  assign n6330 = n3484 & ~n5309 ;
  assign n6331 = ~n6329 & ~n6330 ;
  assign n6332 = ~n3484 & ~n5383 ;
  assign n6333 = n3484 & ~n5396 ;
  assign n6334 = ~n6332 & ~n6333 ;
  assign n6335 = ~n3484 & ~n5470 ;
  assign n6336 = n3484 & ~n5483 ;
  assign n6337 = ~n6335 & ~n6336 ;
  assign n6338 = ~n3484 & ~n5557 ;
  assign n6339 = n3484 & ~n5570 ;
  assign n6340 = ~n6338 & ~n6339 ;
  assign n6341 = ~n3484 & ~n5644 ;
  assign n6342 = n3484 & ~n5657 ;
  assign n6343 = ~n6341 & ~n6342 ;
  assign n6344 = ~n3484 & ~n5731 ;
  assign n6345 = n3484 & ~n5744 ;
  assign n6346 = ~n6344 & ~n6345 ;
  assign n6347 = ~n3484 & ~n5818 ;
  assign n6348 = n3484 & ~n5831 ;
  assign n6349 = ~n6347 & ~n6348 ;
  assign n6350 = ~n3484 & ~n5905 ;
  assign n6351 = n3484 & ~n5918 ;
  assign n6352 = ~n6350 & ~n6351 ;
  assign n6353 = ~n3484 & ~n5992 ;
  assign n6354 = n3484 & ~n6005 ;
  assign n6355 = ~n6353 & ~n6354 ;
  assign n6356 = ~n3484 & ~n6079 ;
  assign n6357 = n3484 & ~n6092 ;
  assign n6358 = ~n6356 & ~n6357 ;
  assign n6359 = ~n3484 & ~n6166 ;
  assign n6360 = n3484 & ~n6179 ;
  assign n6361 = ~n6359 & ~n6360 ;
  assign n6362 = ~n3484 & ~n6253 ;
  assign n6363 = n3484 & ~n6266 ;
  assign n6364 = ~n6362 & ~n6363 ;
  assign n6365 = n3439 & ~n3553 ;
  assign n6366 = ~n3439 & ~n3563 ;
  assign n6367 = ~n6365 & ~n6366 ;
  assign n6368 = ~n3439 & ~n3647 ;
  assign n6369 = n3439 & ~n3654 ;
  assign n6370 = ~n6368 & ~n6369 ;
  assign n6371 = ~n3439 & ~n3734 ;
  assign n6372 = n3439 & ~n3741 ;
  assign n6373 = ~n6371 & ~n6372 ;
  assign n6374 = ~n3439 & ~n3821 ;
  assign n6375 = n3439 & ~n3828 ;
  assign n6376 = ~n6374 & ~n6375 ;
  assign n6377 = ~n3439 & ~n3908 ;
  assign n6378 = n3439 & ~n3915 ;
  assign n6379 = ~n6377 & ~n6378 ;
  assign n6380 = ~n3439 & ~n3995 ;
  assign n6381 = n3439 & ~n4002 ;
  assign n6382 = ~n6380 & ~n6381 ;
  assign n6383 = ~n3439 & ~n4082 ;
  assign n6384 = n3439 & ~n4089 ;
  assign n6385 = ~n6383 & ~n6384 ;
  assign n6386 = ~n3439 & ~n4169 ;
  assign n6387 = n3439 & ~n4176 ;
  assign n6388 = ~n6386 & ~n6387 ;
  assign n6389 = ~n3439 & ~n4256 ;
  assign n6390 = n3439 & ~n4263 ;
  assign n6391 = ~n6389 & ~n6390 ;
  assign n6392 = ~n3439 & ~n4343 ;
  assign n6393 = n3439 & ~n4350 ;
  assign n6394 = ~n6392 & ~n6393 ;
  assign n6395 = ~n3439 & ~n4430 ;
  assign n6396 = n3439 & ~n4437 ;
  assign n6397 = ~n6395 & ~n6396 ;
  assign n6398 = ~n3439 & ~n4517 ;
  assign n6399 = n3439 & ~n4524 ;
  assign n6400 = ~n6398 & ~n6399 ;
  assign n6401 = ~n3439 & ~n4604 ;
  assign n6402 = n3439 & ~n4611 ;
  assign n6403 = ~n6401 & ~n6402 ;
  assign n6404 = ~n3439 & ~n4691 ;
  assign n6405 = n3439 & ~n4698 ;
  assign n6406 = ~n6404 & ~n6405 ;
  assign n6407 = ~n3439 & ~n4778 ;
  assign n6408 = n3439 & ~n4785 ;
  assign n6409 = ~n6407 & ~n6408 ;
  assign n6410 = ~n3439 & ~n4865 ;
  assign n6411 = n3439 & ~n4872 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = ~n3439 & ~n4952 ;
  assign n6414 = n3439 & ~n4959 ;
  assign n6415 = ~n6413 & ~n6414 ;
  assign n6416 = ~n3439 & ~n5039 ;
  assign n6417 = n3439 & ~n5046 ;
  assign n6418 = ~n6416 & ~n6417 ;
  assign n6419 = ~n3439 & ~n5126 ;
  assign n6420 = n3439 & ~n5133 ;
  assign n6421 = ~n6419 & ~n6420 ;
  assign n6422 = ~n3439 & ~n5213 ;
  assign n6423 = n3439 & ~n5220 ;
  assign n6424 = ~n6422 & ~n6423 ;
  assign n6425 = ~n3439 & ~n5300 ;
  assign n6426 = n3439 & ~n5307 ;
  assign n6427 = ~n6425 & ~n6426 ;
  assign n6428 = ~n3439 & ~n5387 ;
  assign n6429 = n3439 & ~n5394 ;
  assign n6430 = ~n6428 & ~n6429 ;
  assign n6431 = ~n3439 & ~n5474 ;
  assign n6432 = n3439 & ~n5481 ;
  assign n6433 = ~n6431 & ~n6432 ;
  assign n6434 = ~n3439 & ~n5561 ;
  assign n6435 = n3439 & ~n5568 ;
  assign n6436 = ~n6434 & ~n6435 ;
  assign n6437 = ~n3439 & ~n5648 ;
  assign n6438 = n3439 & ~n5655 ;
  assign n6439 = ~n6437 & ~n6438 ;
  assign n6440 = ~n3439 & ~n5735 ;
  assign n6441 = n3439 & ~n5742 ;
  assign n6442 = ~n6440 & ~n6441 ;
  assign n6443 = ~n3439 & ~n5822 ;
  assign n6444 = n3439 & ~n5829 ;
  assign n6445 = ~n6443 & ~n6444 ;
  assign n6446 = ~n3439 & ~n5909 ;
  assign n6447 = n3439 & ~n5916 ;
  assign n6448 = ~n6446 & ~n6447 ;
  assign n6449 = ~n3439 & ~n5996 ;
  assign n6450 = n3439 & ~n6003 ;
  assign n6451 = ~n6449 & ~n6450 ;
  assign n6452 = ~n3439 & ~n6083 ;
  assign n6453 = n3439 & ~n6090 ;
  assign n6454 = ~n6452 & ~n6453 ;
  assign n6455 = ~n3439 & ~n6170 ;
  assign n6456 = n3439 & ~n6177 ;
  assign n6457 = ~n6455 & ~n6456 ;
  assign n6458 = ~n3439 & ~n6257 ;
  assign n6459 = n3439 & ~n6264 ;
  assign n6460 = ~n6458 & ~n6459 ;
  assign y0 = ~n3571 ;
  assign y1 = ~n3658 ;
  assign y2 = ~n3745 ;
  assign y3 = ~n3832 ;
  assign y4 = ~n3919 ;
  assign y5 = ~n4006 ;
  assign y6 = ~n4093 ;
  assign y7 = ~n4180 ;
  assign y8 = ~n4267 ;
  assign y9 = ~n4354 ;
  assign y10 = ~n4441 ;
  assign y11 = ~n4528 ;
  assign y12 = ~n4615 ;
  assign y13 = ~n4702 ;
  assign y14 = ~n4789 ;
  assign y15 = ~n4876 ;
  assign y16 = ~n4963 ;
  assign y17 = ~n5050 ;
  assign y18 = ~n5137 ;
  assign y19 = ~n5224 ;
  assign y20 = ~n5311 ;
  assign y21 = ~n5398 ;
  assign y22 = ~n5485 ;
  assign y23 = ~n5572 ;
  assign y24 = ~n5659 ;
  assign y25 = ~n5746 ;
  assign y26 = ~n5833 ;
  assign y27 = ~n5920 ;
  assign y28 = ~n6007 ;
  assign y29 = ~n6094 ;
  assign y30 = ~n6181 ;
  assign y31 = ~n6268 ;
  assign y32 = ~n6271 ;
  assign y33 = ~n6274 ;
  assign y34 = ~n6277 ;
  assign y35 = ~n6280 ;
  assign y36 = ~n6283 ;
  assign y37 = ~n6286 ;
  assign y38 = ~n6289 ;
  assign y39 = ~n6292 ;
  assign y40 = ~n6295 ;
  assign y41 = ~n6298 ;
  assign y42 = ~n6301 ;
  assign y43 = ~n6304 ;
  assign y44 = ~n6307 ;
  assign y45 = ~n6310 ;
  assign y46 = ~n6313 ;
  assign y47 = ~n6316 ;
  assign y48 = ~n6319 ;
  assign y49 = ~n6322 ;
  assign y50 = ~n6325 ;
  assign y51 = ~n6328 ;
  assign y52 = ~n6331 ;
  assign y53 = ~n6334 ;
  assign y54 = ~n6337 ;
  assign y55 = ~n6340 ;
  assign y56 = ~n6343 ;
  assign y57 = ~n6346 ;
  assign y58 = ~n6349 ;
  assign y59 = ~n6352 ;
  assign y60 = ~n6355 ;
  assign y61 = ~n6358 ;
  assign y62 = ~n6361 ;
  assign y63 = ~n6364 ;
  assign y64 = ~n6367 ;
  assign y65 = ~n6370 ;
  assign y66 = ~n6373 ;
  assign y67 = ~n6376 ;
  assign y68 = ~n6379 ;
  assign y69 = ~n6382 ;
  assign y70 = ~n6385 ;
  assign y71 = ~n6388 ;
  assign y72 = ~n6391 ;
  assign y73 = ~n6394 ;
  assign y74 = ~n6397 ;
  assign y75 = ~n6400 ;
  assign y76 = ~n6403 ;
  assign y77 = ~n6406 ;
  assign y78 = ~n6409 ;
  assign y79 = ~n6412 ;
  assign y80 = ~n6415 ;
  assign y81 = ~n6418 ;
  assign y82 = ~n6421 ;
  assign y83 = ~n6424 ;
  assign y84 = ~n6427 ;
  assign y85 = ~n6430 ;
  assign y86 = ~n6433 ;
  assign y87 = ~n6436 ;
  assign y88 = ~n6439 ;
  assign y89 = ~n6442 ;
  assign y90 = ~n6445 ;
  assign y91 = ~n6448 ;
  assign y92 = ~n6451 ;
  assign y93 = ~n6454 ;
  assign y94 = ~n6457 ;
  assign y95 = ~n6460 ;
endmodule
