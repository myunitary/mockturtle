module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 ;
  assign n77 = x9 & x10 ;
  assign n78 = n77 ^ x9 ;
  assign n79 = n78 ^ x10 ;
  assign n259 = n79 ^ x11 ;
  assign n260 = n79 ^ x12 ;
  assign n261 = n259 & n260 ;
  assign n262 = n261 ^ n260 ;
  assign n80 = x11 & x14 ;
  assign n81 = n79 & n80 ;
  assign n70 = x12 & x13 ;
  assign n71 = n70 ^ x12 ;
  assign n72 = n71 ^ x13 ;
  assign n74 = x15 & x16 ;
  assign n264 = ~n72 & n74 ;
  assign n265 = n81 & n264 ;
  assign n73 = x14 & n72 ;
  assign n263 = n73 & n74 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = n266 ^ n74 ;
  assign n268 = n267 ^ n74 ;
  assign n269 = n268 ^ x15 ;
  assign n89 = x11 & n79 ;
  assign n90 = n89 ^ x11 ;
  assign n91 = n90 ^ x11 ;
  assign n85 = n73 ^ x14 ;
  assign n88 = n85 ^ n72 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n89 ^ n72 ;
  assign n94 = n92 & n93 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n97 ^ n92 ;
  assign n86 = n85 ^ x14 ;
  assign n87 = n86 ^ n72 ;
  assign n99 = n98 ^ n87 ;
  assign n100 = n99 ^ n89 ;
  assign n270 = n269 ^ n100 ;
  assign n278 = ~n262 & ~n270 ;
  assign n279 = n278 ^ n270 ;
  assign n280 = n279 ^ n262 ;
  assign n160 = x20 & x21 ;
  assign n161 = n160 ^ x20 ;
  assign n162 = x22 & x23 ;
  assign n163 = n162 ^ x23 ;
  assign n221 = ~x1 & ~x2 ;
  assign n222 = ~n163 & n221 ;
  assign n223 = n222 ^ n221 ;
  assign n224 = ~n161 & n223 ;
  assign n225 = n224 ^ n223 ;
  assign n226 = x24 & x25 ;
  assign n227 = x26 & n226 ;
  assign n228 = n227 ^ n226 ;
  assign n229 = x13 & x14 ;
  assign n230 = n229 ^ x14 ;
  assign n231 = x18 & x19 ;
  assign n232 = n231 ^ x19 ;
  assign n233 = n230 & n232 ;
  assign n234 = n233 ^ n230 ;
  assign n235 = n234 ^ n232 ;
  assign n236 = n235 ^ n230 ;
  assign n237 = n236 ^ n232 ;
  assign n238 = n228 & ~n237 ;
  assign n239 = n238 ^ n228 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n240 ^ n237 ;
  assign n242 = x5 & x6 ;
  assign n243 = n242 ^ x5 ;
  assign n244 = n243 ^ x6 ;
  assign n245 = n78 & n244 ;
  assign n246 = n245 ^ n78 ;
  assign n247 = x3 & x4 ;
  assign n248 = n247 ^ x3 ;
  assign n249 = n248 ^ x4 ;
  assign n250 = x7 & x8 ;
  assign n251 = n250 ^ x7 ;
  assign n252 = n251 ^ x8 ;
  assign n253 = n249 & ~n252 ;
  assign n254 = n253 ^ n252 ;
  assign n255 = n246 & ~n254 ;
  assign n256 = ~n241 & n255 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = n225 & n257 ;
  assign n271 = ~n262 & n270 ;
  assign n272 = n271 ^ n262 ;
  assign n273 = n272 ^ n270 ;
  assign n274 = n258 & n273 ;
  assign n275 = n274 ^ n273 ;
  assign n276 = n275 ^ n258 ;
  assign n277 = n276 ^ n262 ;
  assign n281 = n280 ^ n277 ;
  assign n282 = n281 ^ n258 ;
  assign n75 = n74 ^ x15 ;
  assign n82 = ~n72 & n75 ;
  assign n83 = n81 & n82 ;
  assign n76 = n73 & n75 ;
  assign n84 = n83 ^ n76 ;
  assign n101 = n100 ^ n84 ;
  assign n102 = n101 ^ n75 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n103 ^ n75 ;
  assign n105 = n104 ^ x16 ;
  assign n106 = x17 & n105 ;
  assign n107 = n106 ^ x17 ;
  assign n108 = n107 ^ x17 ;
  assign n61 = ~x21 & ~x22 ;
  assign n62 = x19 & x20 ;
  assign n197 = n61 & n62 ;
  assign n199 = x17 & ~x18 ;
  assign n200 = n197 & n199 ;
  assign n201 = n105 & n200 ;
  assign n198 = x18 & n197 ;
  assign n202 = n201 ^ n198 ;
  assign n203 = n202 ^ n61 ;
  assign n149 = x27 & x28 ;
  assign n150 = x29 & n149 ;
  assign n204 = x23 & x24 ;
  assign n205 = x25 & ~x26 ;
  assign n206 = n204 & n205 ;
  assign n207 = n150 & n206 ;
  assign n208 = ~n203 & n207 ;
  assign n196 = x26 & n150 ;
  assign n209 = n208 ^ n196 ;
  assign n283 = n108 & n209 ;
  assign n284 = ~n282 & n283 ;
  assign n151 = x19 & x25 ;
  assign n152 = x26 & n151 ;
  assign n153 = n152 ^ n151 ;
  assign n154 = n72 & ~n75 ;
  assign n155 = n154 ^ n72 ;
  assign n156 = n155 ^ n75 ;
  assign n157 = ~n153 & n156 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n150 & n158 ;
  assign n164 = ~n161 & ~n163 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = x0 & x1 ;
  assign n168 = n79 & n167 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = ~n166 & ~n169 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = x6 & x7 ;
  assign n173 = x8 & x11 ;
  assign n174 = n172 & n173 ;
  assign n175 = x2 & x3 ;
  assign n176 = x4 & x5 ;
  assign n177 = n175 & n176 ;
  assign n178 = n174 & n177 ;
  assign n179 = ~n171 & n178 ;
  assign n180 = n159 & n179 ;
  assign n181 = n72 & ~n89 ;
  assign n182 = n181 ^ n89 ;
  assign n183 = n182 ^ x14 ;
  assign n184 = n180 & n183 ;
  assign n185 = n184 ^ n180 ;
  assign n186 = n185 ^ n180 ;
  assign n187 = n105 ^ x17 ;
  assign n188 = x18 & n187 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = n186 & n189 ;
  assign n215 = n190 ^ n189 ;
  assign n216 = n215 ^ n189 ;
  assign n217 = n209 & n216 ;
  assign n137 = x23 & ~n61 ;
  assign n138 = ~x23 & n61 ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = x18 & ~n62 ;
  assign n141 = ~x18 & n62 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n139 & ~n142 ;
  assign n144 = ~n139 & n142 ;
  assign n145 = ~n143 & ~n144 ;
  assign n63 = n62 ^ n61 ;
  assign n67 = n61 ^ x18 ;
  assign n68 = n63 & ~n67 ;
  assign n69 = n68 ^ x18 ;
  assign n117 = n69 ^ n62 ;
  assign n118 = n117 ^ n61 ;
  assign n119 = n118 ^ x23 ;
  assign n121 = x17 & n119 ;
  assign n122 = n105 & n121 ;
  assign n120 = ~n69 & n119 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n123 ^ n119 ;
  assign n125 = n124 ^ n69 ;
  assign n126 = n125 ^ n108 ;
  assign n109 = n108 ^ n69 ;
  assign n64 = x23 & ~n63 ;
  assign n65 = ~x23 & n63 ;
  assign n66 = ~n64 & ~n65 ;
  assign n110 = n109 ^ n66 ;
  assign n111 = n108 ^ n62 ;
  assign n112 = n111 ^ n69 ;
  assign n113 = n110 & n112 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ n110 ;
  assign n116 = n115 ^ n112 ;
  assign n127 = n126 ^ n116 ;
  assign n128 = n127 ^ n69 ;
  assign n129 = n128 ^ n66 ;
  assign n130 = n108 ^ x23 ;
  assign n131 = n130 ^ n126 ;
  assign n132 = n129 & n131 ;
  assign n133 = n132 ^ n129 ;
  assign n134 = n133 ^ n116 ;
  assign n135 = n134 ^ n126 ;
  assign n136 = n135 ^ n68 ;
  assign n146 = n145 ^ n136 ;
  assign n147 = n146 ^ x23 ;
  assign n148 = n147 ^ x24 ;
  assign n191 = n190 ^ n148 ;
  assign n210 = n148 & n209 ;
  assign n211 = n210 ^ n209 ;
  assign n212 = n191 & n211 ;
  assign n213 = n212 ^ n211 ;
  assign n214 = n213 ^ n211 ;
  assign n218 = n217 ^ n214 ;
  assign n192 = n148 & n191 ;
  assign n193 = n192 ^ n148 ;
  assign n194 = n193 ^ n191 ;
  assign n195 = n194 ^ n148 ;
  assign n219 = n218 ^ n195 ;
  assign n220 = n219 ^ n216 ;
  assign n285 = n284 ^ n220 ;
  assign n585 = n187 ^ n186 ;
  assign n623 = n585 ^ x18 ;
  assign n333 = x54 & x55 ;
  assign n334 = x30 & x31 ;
  assign n335 = n333 & n334 ;
  assign n317 = x39 & x40 ;
  assign n318 = n317 ^ x39 ;
  assign n319 = n318 ^ x40 ;
  assign n336 = x48 & x49 ;
  assign n337 = n336 ^ x48 ;
  assign n338 = n337 ^ x49 ;
  assign n339 = n319 & ~n338 ;
  assign n340 = n339 ^ n319 ;
  assign n341 = n340 ^ n338 ;
  assign n342 = n335 & ~n341 ;
  assign n343 = n342 ^ n335 ;
  assign n315 = x43 & x44 ;
  assign n316 = n315 ^ x44 ;
  assign n367 = n316 ^ n315 ;
  assign n320 = x41 & x42 ;
  assign n321 = n320 ^ x41 ;
  assign n322 = n319 & n321 ;
  assign n323 = n322 ^ n321 ;
  assign n324 = n323 ^ n321 ;
  assign n325 = n324 ^ x42 ;
  assign n366 = n325 ^ n315 ;
  assign n368 = n367 ^ n366 ;
  assign n394 = n367 ^ n315 ;
  assign n395 = n368 & n394 ;
  assign n396 = n395 ^ n367 ;
  assign n397 = n343 & n396 ;
  assign n398 = n397 ^ n343 ;
  assign n372 = x45 & x46 ;
  assign n373 = n372 ^ x45 ;
  assign n375 = n316 & n373 ;
  assign n376 = n325 & n375 ;
  assign n374 = n315 & n373 ;
  assign n377 = n376 ^ n374 ;
  assign n369 = n366 ^ n315 ;
  assign n370 = n368 & n369 ;
  assign n371 = n370 ^ n366 ;
  assign n378 = n377 ^ n371 ;
  assign n379 = n378 ^ n371 ;
  assign n380 = n379 ^ x46 ;
  assign n399 = x47 & ~x49 ;
  assign n400 = n380 & n399 ;
  assign n401 = ~n398 & n400 ;
  assign n402 = n401 ^ n400 ;
  assign n298 = x36 & x37 ;
  assign n299 = x38 & x41 ;
  assign n300 = n298 & n299 ;
  assign n301 = x32 & x33 ;
  assign n302 = x34 & x35 ;
  assign n303 = n301 & n302 ;
  assign n304 = n300 & n303 ;
  assign n305 = x57 & x58 ;
  assign n306 = x59 & n305 ;
  assign n307 = n304 & n306 ;
  assign n308 = x46 & x47 ;
  assign n309 = n308 ^ x47 ;
  assign n310 = x50 & x56 ;
  assign n311 = n310 ^ x50 ;
  assign n312 = ~n309 & ~n311 ;
  assign n313 = n312 ^ n309 ;
  assign n314 = n313 ^ n311 ;
  assign n358 = ~x43 & x44 ;
  assign n359 = ~n325 & n358 ;
  assign n360 = n359 ^ x44 ;
  assign n361 = n360 ^ x45 ;
  assign n345 = x44 & x45 ;
  assign n346 = n345 ^ x45 ;
  assign n350 = x43 & ~n346 ;
  assign n351 = n350 ^ x43 ;
  assign n352 = n319 & n320 ;
  assign n353 = n352 ^ x43 ;
  assign n354 = ~n351 & n353 ;
  assign n347 = n346 ^ x43 ;
  assign n348 = ~n346 & ~n347 ;
  assign n349 = n348 ^ n346 ;
  assign n355 = n354 ^ n349 ;
  assign n356 = n355 ^ n352 ;
  assign n357 = n356 ^ n346 ;
  assign n362 = n361 ^ n357 ;
  assign n403 = ~n314 & n362 ;
  assign n404 = n403 ^ n314 ;
  assign n405 = n307 & ~n404 ;
  assign n406 = n402 & n405 ;
  assign n381 = x47 & ~x48 ;
  assign n382 = n380 & n381 ;
  assign n383 = n382 ^ x48 ;
  assign n407 = n406 ^ n383 ;
  assign n408 = n407 ^ n362 ;
  assign n326 = ~n316 & n325 ;
  assign n327 = n326 ^ n316 ;
  assign n328 = n327 ^ n325 ;
  assign n329 = n328 ^ x44 ;
  assign n330 = ~n314 & n329 ;
  assign n331 = n330 ^ n314 ;
  assign n332 = n307 & ~n331 ;
  assign n344 = n343 ^ n332 ;
  assign n363 = n362 ^ n343 ;
  assign n389 = n363 ^ n332 ;
  assign n364 = n362 & ~n363 ;
  assign n365 = n364 ^ n343 ;
  assign n384 = n383 ^ n362 ;
  assign n385 = n384 ^ n343 ;
  assign n386 = ~n365 & ~n385 ;
  assign n387 = n386 ^ n364 ;
  assign n388 = n387 ^ n383 ;
  assign n390 = n389 ^ n388 ;
  assign n391 = n344 & n390 ;
  assign n392 = n391 ^ n386 ;
  assign n393 = n392 ^ n364 ;
  assign n409 = n408 ^ n393 ;
  assign n419 = x53 & n333 ;
  assign n446 = n419 ^ x49 ;
  assign n424 = x51 & x52 ;
  assign n425 = n424 ^ x51 ;
  assign n426 = n425 ^ x52 ;
  assign n435 = n426 ^ x50 ;
  assign n436 = n435 ^ x49 ;
  assign n437 = n426 ^ x49 ;
  assign n438 = n436 & n437 ;
  assign n439 = n438 ^ n436 ;
  assign n440 = n439 ^ n437 ;
  assign n441 = n440 ^ x50 ;
  assign n447 = n446 ^ n441 ;
  assign n448 = n447 ^ n381 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = n449 ^ n448 ;
  assign n451 = n450 ^ n381 ;
  assign n452 = n451 ^ n380 ;
  assign n453 = n380 & ~n452 ;
  assign n454 = n453 ^ n452 ;
  assign n455 = n454 ^ n450 ;
  assign n456 = n455 ^ n381 ;
  assign n442 = n441 ^ n419 ;
  assign n443 = n442 ^ x49 ;
  assign n444 = ~x48 & ~n443 ;
  assign n431 = ~x49 & ~x50 ;
  assign n432 = n426 & n431 ;
  assign n433 = n432 ^ x49 ;
  assign n429 = ~x49 & x53 ;
  assign n430 = n333 & n429 ;
  assign n434 = n433 ^ n430 ;
  assign n445 = n444 ^ n434 ;
  assign n457 = n456 ^ n445 ;
  assign n427 = n426 ^ n419 ;
  assign n428 = n419 & ~n427 ;
  assign n458 = n457 ^ n428 ;
  assign n459 = n458 ^ n440 ;
  assign n460 = n459 ^ n436 ;
  assign n420 = x56 & x59 ;
  assign n421 = n420 ^ x59 ;
  assign n422 = n305 & n421 ;
  assign n461 = n419 & n422 ;
  assign n462 = n427 & n461 ;
  assign n463 = n462 ^ n461 ;
  assign n464 = n463 ^ n461 ;
  assign n465 = ~n460 & n464 ;
  assign n466 = n465 ^ n464 ;
  assign n423 = ~n419 & n422 ;
  assign n467 = n466 ^ n423 ;
  assign n468 = n467 ^ n306 ;
  assign n410 = x52 & x53 ;
  assign n411 = n410 ^ x53 ;
  assign n412 = x49 & x50 ;
  assign n413 = n411 & n412 ;
  assign n414 = n413 ^ n412 ;
  assign n415 = n383 & n414 ;
  assign n416 = n415 ^ n414 ;
  assign n417 = n416 ^ n414 ;
  assign n418 = n417 ^ n411 ;
  assign n506 = n468 ^ n418 ;
  assign n508 = n414 ^ n411 ;
  assign n509 = n508 ^ n414 ;
  assign n479 = x52 & ~x53 ;
  assign n480 = n412 & ~n479 ;
  assign n507 = n480 ^ n414 ;
  assign n510 = n509 ^ n507 ;
  assign n511 = n507 ^ n414 ;
  assign n512 = ~n510 & n511 ;
  assign n513 = n512 ^ n507 ;
  assign n514 = n383 & n513 ;
  assign n515 = n514 ^ n508 ;
  assign n516 = n515 ^ n414 ;
  assign n517 = n506 & n516 ;
  assign n518 = n517 ^ n516 ;
  assign n485 = n383 & n480 ;
  assign n486 = n485 ^ n480 ;
  assign n487 = n486 ^ n480 ;
  assign n496 = n487 ^ n418 ;
  assign n505 = n487 & n496 ;
  assign n519 = n518 ^ n505 ;
  assign n520 = n519 ^ n468 ;
  assign n521 = n520 ^ n409 ;
  assign n503 = n468 & n487 ;
  assign n504 = n503 ^ n468 ;
  assign n522 = n521 ^ n504 ;
  assign n523 = n409 & n522 ;
  assign n524 = n523 ^ n409 ;
  assign n525 = n524 ^ n522 ;
  assign n526 = n525 ^ n409 ;
  assign n527 = n526 ^ n409 ;
  assign n528 = n527 ^ n522 ;
  assign n495 = n487 ^ n468 ;
  assign n497 = ~n418 & n496 ;
  assign n498 = n497 ^ n418 ;
  assign n499 = n498 ^ n468 ;
  assign n500 = ~n495 & ~n499 ;
  assign n501 = n500 ^ n497 ;
  assign n502 = n501 ^ n468 ;
  assign n529 = n528 ^ n502 ;
  assign n530 = n529 ^ n418 ;
  assign n531 = n530 ^ n468 ;
  assign n532 = x56 & x57 ;
  assign n533 = n532 ^ x57 ;
  assign n534 = x46 & x51 ;
  assign n535 = n534 ^ x46 ;
  assign n536 = n535 ^ x51 ;
  assign n537 = n533 & n536 ;
  assign n538 = n537 ^ n533 ;
  assign n539 = x41 & x43 ;
  assign n540 = n539 ^ x41 ;
  assign n541 = n345 & n540 ;
  assign n542 = n538 & n541 ;
  assign n543 = x37 & x38 ;
  assign n544 = n543 ^ x37 ;
  assign n545 = n544 ^ x38 ;
  assign n546 = n318 & n545 ;
  assign n547 = n546 ^ n318 ;
  assign n548 = x41 & n319 ;
  assign n549 = n548 ^ x42 ;
  assign n550 = n547 & n549 ;
  assign n551 = n542 & n550 ;
  assign n552 = x47 & x48 ;
  assign n553 = n414 ^ n412 ;
  assign n554 = n552 & n553 ;
  assign n555 = n554 ^ n553 ;
  assign n556 = x33 & x34 ;
  assign n557 = n556 ^ x33 ;
  assign n558 = n557 ^ x34 ;
  assign n559 = x35 & x36 ;
  assign n560 = n559 ^ x35 ;
  assign n561 = n560 ^ x36 ;
  assign n562 = n558 & n561 ;
  assign n563 = n562 ^ n558 ;
  assign n564 = n563 ^ n561 ;
  assign n565 = x31 & x32 ;
  assign n566 = n565 ^ x31 ;
  assign n567 = n566 ^ x32 ;
  assign n568 = n333 & n567 ;
  assign n569 = n568 ^ n333 ;
  assign n570 = ~n564 & n569 ;
  assign n571 = n555 & n570 ;
  assign n572 = n551 & n571 ;
  assign n573 = ~x0 & ~x30 ;
  assign n608 = x48 ^ x47 ;
  assign n609 = n380 & n608 ;
  assign n610 = n609 ^ x48 ;
  assign n613 = n573 & n610 ;
  assign n614 = n572 & n613 ;
  assign n615 = ~n531 & n614 ;
  assign n616 = n615 ^ n614 ;
  assign n617 = n616 ^ n531 ;
  assign n611 = n572 & n610 ;
  assign n612 = n573 & n611 ;
  assign n618 = n617 ^ n612 ;
  assign n474 = n380 ^ x48 ;
  assign n473 = n381 ^ x48 ;
  assign n475 = n474 ^ n473 ;
  assign n476 = n474 ^ x48 ;
  assign n477 = n475 & n476 ;
  assign n478 = n477 ^ n474 ;
  assign n469 = ~x0 & ~x51 ;
  assign n481 = ~n469 & n480 ;
  assign n482 = n478 & n481 ;
  assign n483 = n468 & n482 ;
  assign n484 = n483 ^ n482 ;
  assign n488 = n487 ^ n484 ;
  assign n470 = n468 & n469 ;
  assign n471 = n470 ^ n468 ;
  assign n472 = n471 ^ n469 ;
  assign n489 = n488 ^ n472 ;
  assign n597 = n409 & n418 ;
  assign n598 = n597 ^ n409 ;
  assign n599 = n598 ^ n418 ;
  assign n600 = n599 ^ n418 ;
  assign n601 = n600 ^ n409 ;
  assign n602 = n601 ^ n418 ;
  assign n603 = n489 & ~n602 ;
  assign n604 = n603 ^ n489 ;
  assign n605 = n604 ^ n602 ;
  assign n606 = n605 ^ n489 ;
  assign n607 = n606 ^ n602 ;
  assign n619 = n618 ^ n607 ;
  assign n620 = n619 ^ n489 ;
  assign n592 = n189 ^ n148 ;
  assign n621 = n620 ^ n592 ;
  assign n586 = x18 & ~n187 ;
  assign n587 = n586 ^ n186 ;
  assign n588 = n587 ^ x18 ;
  assign n589 = n585 & ~n588 ;
  assign n590 = n589 ^ n586 ;
  assign n584 = n187 ^ x18 ;
  assign n591 = n590 ^ n584 ;
  assign n593 = n592 ^ n589 ;
  assign n594 = n593 ^ n186 ;
  assign n595 = ~n591 & ~n594 ;
  assign n596 = n595 ^ n586 ;
  assign n622 = n621 ^ n596 ;
  assign n624 = n623 ^ n622 ;
  assign n292 = ~n108 & n282 ;
  assign n293 = n292 ^ n108 ;
  assign n294 = n293 ^ n282 ;
  assign n625 = n624 ^ n294 ;
  assign n628 = n108 & ~n209 ;
  assign n629 = ~n282 & n628 ;
  assign n286 = ~x18 & n183 ;
  assign n287 = n187 & n286 ;
  assign n288 = n180 & n287 ;
  assign n289 = n148 & n288 ;
  assign n290 = n289 ^ n288 ;
  assign n291 = n290 ^ n216 ;
  assign n626 = n209 & n291 ;
  assign n627 = n626 ^ n291 ;
  assign n630 = n629 ^ n627 ;
  assign n631 = n625 & n630 ;
  assign n632 = n631 ^ n630 ;
  assign n633 = n632 ^ n630 ;
  assign n634 = n633 ^ n630 ;
  assign n575 = x47 & n380 ;
  assign n576 = x48 & ~n380 ;
  assign n577 = n573 & ~n576 ;
  assign n578 = ~n575 & n577 ;
  assign n579 = n572 & n578 ;
  assign n574 = n572 & n573 ;
  assign n580 = n579 ^ n574 ;
  assign n581 = n294 & ~n580 ;
  assign n582 = ~n531 & n581 ;
  assign n295 = n294 ^ n291 ;
  assign n296 = n295 ^ n291 ;
  assign n490 = n418 & n489 ;
  assign n491 = n409 & n490 ;
  assign n492 = n491 ^ n490 ;
  assign n493 = n296 & n492 ;
  assign n494 = n493 ^ n296 ;
  assign n583 = n582 ^ n494 ;
  assign n635 = n634 ^ n583 ;
  assign n297 = ~n209 & n296 ;
  assign n636 = n635 ^ n297 ;
  assign n637 = n636 ^ n620 ;
  assign n638 = n637 ^ n209 ;
  assign n639 = n638 ^ n620 ;
  assign n641 = n284 ^ n209 ;
  assign n640 = n220 ^ n209 ;
  assign n642 = n641 ^ n640 ;
  assign n658 = n262 & ~n270 ;
  assign n659 = n108 & n658 ;
  assign n660 = n258 & n659 ;
  assign n661 = n660 ^ n108 ;
  assign n662 = n661 ^ n108 ;
  assign n663 = n662 ^ n108 ;
  assign n664 = n663 ^ n108 ;
  assign n688 = ~n209 & n664 ;
  assign n689 = n688 ^ n209 ;
  assign n690 = n689 ^ n664 ;
  assign n670 = n203 & n206 ;
  assign n671 = n670 ^ n206 ;
  assign n672 = n671 ^ x26 ;
  assign n673 = n150 & ~n672 ;
  assign n674 = n673 ^ n150 ;
  assign n680 = n664 & ~n674 ;
  assign n679 = n209 & ~n674 ;
  assign n681 = n680 ^ n679 ;
  assign n649 = n611 ^ n572 ;
  assign n650 = n649 ^ n572 ;
  assign n643 = x0 & x30 ;
  assign n644 = n643 ^ n468 ;
  assign n645 = n468 & n644 ;
  assign n646 = n645 ^ n468 ;
  assign n647 = n646 ^ n644 ;
  assign n651 = n650 ^ n647 ;
  assign n652 = n650 ^ n643 ;
  assign n653 = n651 & n652 ;
  assign n654 = n653 ^ n652 ;
  assign n655 = n654 ^ n651 ;
  assign n648 = n647 ^ n468 ;
  assign n656 = n655 ^ n648 ;
  assign n657 = n656 ^ n650 ;
  assign n677 = n209 & ~n664 ;
  assign n678 = ~n657 & n677 ;
  assign n682 = n681 ^ n678 ;
  assign n676 = n664 ^ n209 ;
  assign n683 = n682 ^ n676 ;
  assign n665 = n664 ^ n657 ;
  assign n666 = n657 & n665 ;
  assign n668 = n666 ^ n657 ;
  assign n669 = n668 ^ n665 ;
  assign n675 = n674 ^ n669 ;
  assign n684 = n683 ^ n675 ;
  assign n667 = n666 ^ n665 ;
  assign n685 = n684 ^ n667 ;
  assign n686 = n685 ^ n674 ;
  assign n687 = n686 ^ n641 ;
  assign n691 = n690 ^ n687 ;
  assign n692 = n642 & n691 ;
  assign n693 = n692 ^ n691 ;
  assign n694 = n693 ^ n691 ;
  assign n695 = n694 ^ n691 ;
  assign n696 = n695 ^ n691 ;
  assign n697 = n696 ^ n642 ;
  assign n698 = n697 ^ n691 ;
  assign n699 = n698 ^ n687 ;
  assign n700 = n699 ^ n640 ;
  assign y0 = ~n285 ;
  assign y1 = ~n639 ;
  assign y2 = n700 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
