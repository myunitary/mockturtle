module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n9 = x6 & x7 ;
  assign n10 = x4 & x5 ;
  assign n11 = n9 & n10 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n12 ^ n10 ;
  assign n27 = x1 & x2 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = x3 & n28 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = ~n13 & n30 ;
  assign n14 = x0 & x1 ;
  assign n23 = n14 ^ x0 ;
  assign n24 = x3 & n23 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~n13 & n25 ;
  assign n32 = n31 ^ n26 ;
  assign n20 = ~x0 & ~x2 ;
  assign n21 = ~n13 & n20 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = x2 & x3 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = n15 & n17 ;
  assign n19 = ~n13 & n18 ;
  assign n22 = n21 ^ n19 ;
  assign n33 = n32 ^ n22 ;
  assign n42 = n10 ^ x4 ;
  assign n43 = n42 ^ x5 ;
  assign n50 = n33 & ~n43 ;
  assign n34 = n23 ^ x1 ;
  assign n35 = n16 ^ x2 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = ~n34 & ~n36 ;
  assign n38 = n9 ^ x6 ;
  assign n39 = n38 ^ x7 ;
  assign n44 = ~n39 & ~n43 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n37 & ~n45 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n33 & ~n47 ;
  assign n40 = n37 & ~n39 ;
  assign n41 = n33 & n40 ;
  assign n49 = n48 ^ n41 ;
  assign n51 = n50 ^ n49 ;
  assign y0 = n51 ;
endmodule
