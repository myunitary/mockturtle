module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 ;
  assign n168 = x32 ^ x0 ;
  assign n212 = x31 & ~x63 ;
  assign n137 = x63 ^ x31 ;
  assign n210 = x30 & ~x62 ;
  assign n211 = ~n137 & n210 ;
  assign n213 = n212 ^ n211 ;
  assign n138 = x62 ^ x30 ;
  assign n139 = ~n137 & ~n138 ;
  assign n207 = x29 & ~x61 ;
  assign n140 = x61 ^ x29 ;
  assign n205 = x28 & ~x60 ;
  assign n206 = ~n140 & n205 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = n139 & n208 ;
  assign n214 = n213 ^ n209 ;
  assign n141 = x60 ^ x28 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n139 & n142 ;
  assign n201 = x27 & ~x59 ;
  assign n144 = x59 ^ x27 ;
  assign n199 = x26 & ~x58 ;
  assign n200 = ~n144 & n199 ;
  assign n202 = n201 ^ n200 ;
  assign n145 = x58 ^ x26 ;
  assign n146 = ~n144 & ~n145 ;
  assign n196 = x25 & ~x57 ;
  assign n147 = x57 ^ x25 ;
  assign n194 = x24 & ~x56 ;
  assign n195 = ~n147 & n194 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n146 & n197 ;
  assign n203 = n202 ^ n198 ;
  assign n204 = n143 & n203 ;
  assign n215 = n214 ^ n204 ;
  assign n148 = x56 ^ x24 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n146 & n149 ;
  assign n151 = n143 & n150 ;
  assign n189 = x23 & ~x55 ;
  assign n152 = x55 ^ x23 ;
  assign n187 = x22 & ~x54 ;
  assign n188 = ~n152 & n187 ;
  assign n190 = n189 ^ n188 ;
  assign n153 = x54 ^ x22 ;
  assign n154 = ~n152 & ~n153 ;
  assign n184 = x21 & ~x53 ;
  assign n155 = x53 ^ x21 ;
  assign n182 = x20 & ~x52 ;
  assign n183 = ~n155 & n182 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = n154 & n185 ;
  assign n191 = n190 ^ n186 ;
  assign n156 = x52 ^ x20 ;
  assign n157 = ~n155 & ~n156 ;
  assign n158 = n154 & n157 ;
  assign n178 = x19 & ~x51 ;
  assign n159 = x51 ^ x19 ;
  assign n176 = x18 & ~x50 ;
  assign n177 = ~n159 & n176 ;
  assign n179 = n178 ^ n177 ;
  assign n160 = x50 ^ x18 ;
  assign n161 = ~n159 & ~n160 ;
  assign n173 = x17 & ~x49 ;
  assign n162 = x49 ^ x17 ;
  assign n171 = x16 & ~x48 ;
  assign n172 = ~n162 & n171 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = n161 & n174 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n158 & n180 ;
  assign n192 = n191 ^ n181 ;
  assign n193 = n151 & n192 ;
  assign n216 = n215 ^ n193 ;
  assign n217 = n168 & n216 ;
  assign n132 = x15 & ~x47 ;
  assign n98 = x47 ^ x15 ;
  assign n130 = x14 & ~x46 ;
  assign n131 = ~n98 & n130 ;
  assign n133 = n132 ^ n131 ;
  assign n99 = x46 ^ x14 ;
  assign n100 = ~n98 & ~n99 ;
  assign n127 = x13 & ~x45 ;
  assign n101 = x45 ^ x13 ;
  assign n125 = x12 & ~x44 ;
  assign n126 = ~n101 & n125 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n100 & n128 ;
  assign n134 = n133 ^ n129 ;
  assign n102 = x44 ^ x12 ;
  assign n103 = ~n101 & ~n102 ;
  assign n104 = n100 & n103 ;
  assign n121 = x11 & ~x43 ;
  assign n105 = x43 ^ x11 ;
  assign n119 = x10 & ~x42 ;
  assign n120 = ~n105 & n119 ;
  assign n122 = n121 ^ n120 ;
  assign n106 = x42 ^ x10 ;
  assign n107 = ~n105 & ~n106 ;
  assign n116 = x9 & ~x41 ;
  assign n108 = x41 ^ x9 ;
  assign n114 = x8 & ~x40 ;
  assign n115 = ~n108 & n114 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n107 & n117 ;
  assign n123 = n122 ^ n118 ;
  assign n124 = n104 & n123 ;
  assign n135 = n134 ^ n124 ;
  assign n94 = x7 & ~x39 ;
  assign n79 = x39 ^ x7 ;
  assign n92 = x6 & ~x38 ;
  assign n93 = ~n79 & n92 ;
  assign n95 = n94 ^ n93 ;
  assign n80 = x38 ^ x6 ;
  assign n81 = ~n79 & ~n80 ;
  assign n89 = x5 & ~x37 ;
  assign n82 = x37 ^ x5 ;
  assign n87 = x4 & ~x36 ;
  assign n88 = ~n82 & n87 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n81 & n90 ;
  assign n96 = n95 ^ n91 ;
  assign n76 = x3 & ~x35 ;
  assign n70 = x35 ^ x3 ;
  assign n74 = x2 & ~x34 ;
  assign n75 = ~n70 & n74 ;
  assign n77 = n76 ^ n75 ;
  assign n68 = x1 & ~x33 ;
  assign n65 = x33 ^ x1 ;
  assign n66 = x0 & ~x32 ;
  assign n67 = ~n65 & n66 ;
  assign n69 = n68 ^ n67 ;
  assign n71 = x34 ^ x2 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = n69 & n72 ;
  assign n78 = n77 ^ n73 ;
  assign n83 = x36 ^ x4 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = n81 & n84 ;
  assign n86 = n78 & n85 ;
  assign n97 = n96 ^ n86 ;
  assign n109 = x40 ^ x8 ;
  assign n110 = ~n108 & ~n109 ;
  assign n111 = n107 & n110 ;
  assign n112 = n104 & n111 ;
  assign n113 = n97 & n112 ;
  assign n136 = n135 ^ n113 ;
  assign n163 = x48 ^ x16 ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = n161 & n164 ;
  assign n166 = n158 & n165 ;
  assign n167 = n151 & n166 ;
  assign n169 = n167 & n168 ;
  assign n170 = n136 & n169 ;
  assign n218 = n217 ^ n170 ;
  assign n219 = n218 ^ x32 ;
  assign n222 = n65 & n216 ;
  assign n220 = n65 & n167 ;
  assign n221 = n136 & n220 ;
  assign n223 = n222 ^ n221 ;
  assign n224 = n223 ^ x33 ;
  assign n227 = n71 & n216 ;
  assign n225 = n71 & n167 ;
  assign n226 = n136 & n225 ;
  assign n228 = n227 ^ n226 ;
  assign n229 = n228 ^ x34 ;
  assign n232 = n70 & n216 ;
  assign n230 = n70 & n167 ;
  assign n231 = n136 & n230 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = n233 ^ x35 ;
  assign n237 = n83 & n216 ;
  assign n235 = n83 & n167 ;
  assign n236 = n136 & n235 ;
  assign n238 = n237 ^ n236 ;
  assign n239 = n238 ^ x36 ;
  assign n242 = n82 & n216 ;
  assign n240 = n82 & n167 ;
  assign n241 = n136 & n240 ;
  assign n243 = n242 ^ n241 ;
  assign n244 = n243 ^ x37 ;
  assign n247 = n80 & n216 ;
  assign n245 = n80 & n167 ;
  assign n246 = n136 & n245 ;
  assign n248 = n247 ^ n246 ;
  assign n249 = n248 ^ x38 ;
  assign n252 = n79 & n216 ;
  assign n250 = n79 & n167 ;
  assign n251 = n136 & n250 ;
  assign n253 = n252 ^ n251 ;
  assign n254 = n253 ^ x39 ;
  assign n257 = n109 & n216 ;
  assign n255 = n109 & n167 ;
  assign n256 = n136 & n255 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n258 ^ x40 ;
  assign n262 = n108 & n216 ;
  assign n260 = n108 & n167 ;
  assign n261 = n136 & n260 ;
  assign n263 = n262 ^ n261 ;
  assign n264 = n263 ^ x41 ;
  assign n267 = n106 & n216 ;
  assign n265 = n106 & n167 ;
  assign n266 = n136 & n265 ;
  assign n268 = n267 ^ n266 ;
  assign n269 = n268 ^ x42 ;
  assign n272 = n105 & n216 ;
  assign n270 = n105 & n167 ;
  assign n271 = n136 & n270 ;
  assign n273 = n272 ^ n271 ;
  assign n274 = n273 ^ x43 ;
  assign n277 = n102 & n216 ;
  assign n275 = n102 & n167 ;
  assign n276 = n136 & n275 ;
  assign n278 = n277 ^ n276 ;
  assign n279 = n278 ^ x44 ;
  assign n282 = n101 & n216 ;
  assign n280 = n101 & n167 ;
  assign n281 = n136 & n280 ;
  assign n283 = n282 ^ n281 ;
  assign n284 = n283 ^ x45 ;
  assign n287 = n99 & n216 ;
  assign n285 = n99 & n167 ;
  assign n286 = n136 & n285 ;
  assign n288 = n287 ^ n286 ;
  assign n289 = n288 ^ x46 ;
  assign n292 = n98 & n216 ;
  assign n290 = n98 & n167 ;
  assign n291 = n136 & n290 ;
  assign n293 = n292 ^ n291 ;
  assign n294 = n293 ^ x47 ;
  assign n297 = n163 & n216 ;
  assign n295 = n163 & n167 ;
  assign n296 = n136 & n295 ;
  assign n298 = n297 ^ n296 ;
  assign n299 = n298 ^ x48 ;
  assign n302 = n162 & n216 ;
  assign n300 = n162 & n167 ;
  assign n301 = n136 & n300 ;
  assign n303 = n302 ^ n301 ;
  assign n304 = n303 ^ x49 ;
  assign n307 = n160 & n216 ;
  assign n305 = n160 & n167 ;
  assign n306 = n136 & n305 ;
  assign n308 = n307 ^ n306 ;
  assign n309 = n308 ^ x50 ;
  assign n312 = n159 & n216 ;
  assign n310 = n159 & n167 ;
  assign n311 = n136 & n310 ;
  assign n313 = n312 ^ n311 ;
  assign n314 = n313 ^ x51 ;
  assign n317 = n156 & n216 ;
  assign n315 = n156 & n167 ;
  assign n316 = n136 & n315 ;
  assign n318 = n317 ^ n316 ;
  assign n319 = n318 ^ x52 ;
  assign n322 = n155 & n216 ;
  assign n320 = n155 & n167 ;
  assign n321 = n136 & n320 ;
  assign n323 = n322 ^ n321 ;
  assign n324 = n323 ^ x53 ;
  assign n327 = n153 & n216 ;
  assign n325 = n153 & n167 ;
  assign n326 = n136 & n325 ;
  assign n328 = n327 ^ n326 ;
  assign n329 = n328 ^ x54 ;
  assign n332 = n152 & n216 ;
  assign n330 = n152 & n167 ;
  assign n331 = n136 & n330 ;
  assign n333 = n332 ^ n331 ;
  assign n334 = n333 ^ x55 ;
  assign n337 = n148 & n216 ;
  assign n335 = n148 & n167 ;
  assign n336 = n136 & n335 ;
  assign n338 = n337 ^ n336 ;
  assign n339 = n338 ^ x56 ;
  assign n342 = n147 & n216 ;
  assign n340 = n147 & n167 ;
  assign n341 = n136 & n340 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = n343 ^ x57 ;
  assign n347 = n145 & n216 ;
  assign n345 = n145 & n167 ;
  assign n346 = n136 & n345 ;
  assign n348 = n347 ^ n346 ;
  assign n349 = n348 ^ x58 ;
  assign n352 = n144 & n216 ;
  assign n350 = n144 & n167 ;
  assign n351 = n136 & n350 ;
  assign n353 = n352 ^ n351 ;
  assign n354 = n353 ^ x59 ;
  assign n357 = n141 & n216 ;
  assign n355 = n141 & n167 ;
  assign n356 = n136 & n355 ;
  assign n358 = n357 ^ n356 ;
  assign n359 = n358 ^ x60 ;
  assign n362 = n140 & n216 ;
  assign n360 = n140 & n167 ;
  assign n361 = n136 & n360 ;
  assign n363 = n362 ^ n361 ;
  assign n364 = n363 ^ x61 ;
  assign n367 = n138 & n216 ;
  assign n365 = n138 & n167 ;
  assign n366 = n136 & n365 ;
  assign n368 = n367 ^ n366 ;
  assign n369 = n368 ^ x62 ;
  assign n372 = n137 & n216 ;
  assign n370 = n137 & n167 ;
  assign n371 = n136 & n370 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = n373 ^ x63 ;
  assign y0 = n219 ;
  assign y1 = n224 ;
  assign y2 = n229 ;
  assign y3 = n234 ;
  assign y4 = n239 ;
  assign y5 = n244 ;
  assign y6 = n249 ;
  assign y7 = n254 ;
  assign y8 = n259 ;
  assign y9 = n264 ;
  assign y10 = n269 ;
  assign y11 = n274 ;
  assign y12 = n279 ;
  assign y13 = n284 ;
  assign y14 = n289 ;
  assign y15 = n294 ;
  assign y16 = n299 ;
  assign y17 = n304 ;
  assign y18 = n309 ;
  assign y19 = n314 ;
  assign y20 = n319 ;
  assign y21 = n324 ;
  assign y22 = n329 ;
  assign y23 = n334 ;
  assign y24 = n339 ;
  assign y25 = n344 ;
  assign y26 = n349 ;
  assign y27 = n354 ;
  assign y28 = n359 ;
  assign y29 = n364 ;
  assign y30 = n369 ;
  assign y31 = n374 ;
endmodule
