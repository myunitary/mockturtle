module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 ;
  assign n73 = x10 ^ x2 ;
  assign n103 = x3 & x11 ;
  assign n104 = n103 ^ x3 ;
  assign n105 = n73 & n104 ;
  assign n106 = n105 ^ n104 ;
  assign n102 = x2 & ~x10 ;
  assign n107 = n106 ^ n102 ;
  assign n68 = x8 ^ x0 ;
  assign n69 = x9 ^ x1 ;
  assign n70 = n68 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n69 ;
  assign n304 = x2 & ~n72 ;
  assign n305 = n107 & n304 ;
  assign n98 = x1 & ~x9 ;
  assign n99 = ~n68 & n98 ;
  assign n97 = x0 & ~x8 ;
  assign n100 = n99 ^ n97 ;
  assign n303 = x2 & ~n100 ;
  assign n306 = n305 ^ n303 ;
  assign n74 = x11 ^ x3 ;
  assign n75 = n73 & n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n72 & n77 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = n79 ^ n77 ;
  assign n50 = x12 ^ x4 ;
  assign n54 = x13 ^ x5 ;
  assign n55 = n50 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = n56 ^ n54 ;
  assign n59 = x14 ^ x6 ;
  assign n84 = x15 ^ x7 ;
  assign n85 = n59 & n84 ;
  assign n86 = n85 ^ n59 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = n57 & n87 ;
  assign n89 = n88 ^ n57 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n80 & n90 ;
  assign n92 = n91 ^ n80 ;
  assign n93 = n92 ^ n90 ;
  assign n300 = x2 & n93 ;
  assign n301 = n300 ^ x2 ;
  assign n302 = n301 ^ x2 ;
  assign n307 = n306 ^ n302 ;
  assign n60 = x7 & x15 ;
  assign n61 = n60 ^ x7 ;
  assign n62 = n59 & n61 ;
  assign n63 = n62 ^ n61 ;
  assign n58 = x6 & ~x14 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = n57 & n64 ;
  assign n66 = n65 ^ n64 ;
  assign n51 = x5 & ~x13 ;
  assign n52 = ~n50 & n51 ;
  assign n49 = x4 & ~x12 ;
  assign n53 = n52 ^ n49 ;
  assign n67 = n66 ^ n53 ;
  assign n297 = x2 & n80 ;
  assign n298 = n297 ^ x2 ;
  assign n299 = n67 & n298 ;
  assign n308 = n307 ^ n299 ;
  assign n291 = x10 & ~n72 ;
  assign n292 = n107 & n291 ;
  assign n290 = x10 & ~n100 ;
  assign n293 = n292 ^ n290 ;
  assign n287 = x10 & n93 ;
  assign n288 = n287 ^ x10 ;
  assign n289 = n288 ^ x10 ;
  assign n294 = n293 ^ n289 ;
  assign n284 = x10 & n80 ;
  assign n285 = n284 ^ x10 ;
  assign n286 = n67 & n285 ;
  assign n295 = n294 ^ n286 ;
  assign n296 = n295 ^ x10 ;
  assign n309 = n308 ^ n296 ;
  assign n310 = n309 ^ x18 ;
  assign n331 = x3 & ~n72 ;
  assign n332 = n107 & n331 ;
  assign n330 = x3 & ~n100 ;
  assign n333 = n332 ^ n330 ;
  assign n327 = x3 & n93 ;
  assign n328 = n327 ^ x3 ;
  assign n329 = n328 ^ x3 ;
  assign n334 = n333 ^ n329 ;
  assign n324 = x3 & n80 ;
  assign n325 = n324 ^ x3 ;
  assign n326 = n67 & n325 ;
  assign n335 = n334 ^ n326 ;
  assign n318 = x11 & ~n72 ;
  assign n319 = n107 & n318 ;
  assign n317 = x11 & ~n100 ;
  assign n320 = n319 ^ n317 ;
  assign n314 = x11 & n93 ;
  assign n315 = n314 ^ x11 ;
  assign n316 = n315 ^ x11 ;
  assign n321 = n320 ^ n316 ;
  assign n311 = x11 & n80 ;
  assign n312 = n311 ^ x11 ;
  assign n313 = n67 & n312 ;
  assign n322 = n321 ^ n313 ;
  assign n323 = n322 ^ x11 ;
  assign n336 = n335 ^ n323 ;
  assign n366 = x19 & n336 ;
  assign n367 = n366 ^ n336 ;
  assign n368 = n310 & n367 ;
  assign n369 = n368 ^ n367 ;
  assign n365 = ~x18 & n309 ;
  assign n370 = n369 ^ n365 ;
  assign n247 = x0 & ~n72 ;
  assign n248 = n107 & n247 ;
  assign n246 = x0 & ~n100 ;
  assign n249 = n248 ^ n246 ;
  assign n243 = x0 & n93 ;
  assign n244 = n243 ^ x0 ;
  assign n245 = n244 ^ x0 ;
  assign n250 = n249 ^ n245 ;
  assign n240 = x0 & n80 ;
  assign n241 = n240 ^ x0 ;
  assign n242 = n67 & n241 ;
  assign n251 = n250 ^ n242 ;
  assign n234 = x8 & ~n72 ;
  assign n235 = n107 & n234 ;
  assign n233 = x8 & ~n100 ;
  assign n236 = n235 ^ n233 ;
  assign n230 = x8 & n93 ;
  assign n231 = n230 ^ x8 ;
  assign n232 = n231 ^ x8 ;
  assign n237 = n236 ^ n232 ;
  assign n227 = x8 & n80 ;
  assign n228 = n227 ^ x8 ;
  assign n229 = n67 & n228 ;
  assign n238 = n237 ^ n229 ;
  assign n239 = n238 ^ x8 ;
  assign n252 = n251 ^ n239 ;
  assign n253 = n252 ^ x16 ;
  assign n274 = x1 & ~n72 ;
  assign n275 = n107 & n274 ;
  assign n273 = x1 & ~n100 ;
  assign n276 = n275 ^ n273 ;
  assign n270 = x1 & n93 ;
  assign n271 = n270 ^ x1 ;
  assign n272 = n271 ^ x1 ;
  assign n277 = n276 ^ n272 ;
  assign n267 = x1 & n80 ;
  assign n268 = n267 ^ x1 ;
  assign n269 = n67 & n268 ;
  assign n278 = n277 ^ n269 ;
  assign n261 = x9 & ~n72 ;
  assign n262 = n107 & n261 ;
  assign n260 = x9 & ~n100 ;
  assign n263 = n262 ^ n260 ;
  assign n257 = x9 & n93 ;
  assign n258 = n257 ^ x9 ;
  assign n259 = n258 ^ x9 ;
  assign n264 = n263 ^ n259 ;
  assign n254 = x9 & n80 ;
  assign n255 = n254 ^ x9 ;
  assign n256 = n67 & n255 ;
  assign n265 = n264 ^ n256 ;
  assign n266 = n265 ^ x9 ;
  assign n279 = n278 ^ n266 ;
  assign n280 = n279 ^ x17 ;
  assign n281 = n253 & n280 ;
  assign n282 = n281 ^ n253 ;
  assign n283 = n282 ^ n280 ;
  assign n417 = x16 & ~n283 ;
  assign n418 = n370 & n417 ;
  assign n361 = ~x17 & n279 ;
  assign n362 = ~n253 & n361 ;
  assign n360 = ~x16 & n252 ;
  assign n363 = n362 ^ n360 ;
  assign n416 = x16 & ~n363 ;
  assign n419 = n418 ^ n416 ;
  assign n337 = n336 ^ x19 ;
  assign n338 = n310 & n337 ;
  assign n339 = n338 ^ n310 ;
  assign n340 = n339 ^ n337 ;
  assign n341 = n283 & n340 ;
  assign n342 = n341 ^ n283 ;
  assign n343 = n342 ^ n340 ;
  assign n121 = x4 & ~n72 ;
  assign n122 = n107 & n121 ;
  assign n120 = x4 & ~n100 ;
  assign n123 = n122 ^ n120 ;
  assign n117 = x4 & n93 ;
  assign n118 = n117 ^ x4 ;
  assign n119 = n118 ^ x4 ;
  assign n124 = n123 ^ n119 ;
  assign n114 = x4 & n80 ;
  assign n115 = n114 ^ x4 ;
  assign n116 = n67 & n115 ;
  assign n125 = n124 ^ n116 ;
  assign n108 = x12 & ~n72 ;
  assign n109 = n107 & n108 ;
  assign n101 = x12 & ~n100 ;
  assign n110 = n109 ^ n101 ;
  assign n94 = x12 & n93 ;
  assign n95 = n94 ^ x12 ;
  assign n96 = n95 ^ x12 ;
  assign n111 = n110 ^ n96 ;
  assign n81 = x12 & n80 ;
  assign n82 = n81 ^ x12 ;
  assign n83 = n67 & n82 ;
  assign n112 = n111 ^ n83 ;
  assign n113 = n112 ^ x12 ;
  assign n126 = n125 ^ n113 ;
  assign n128 = n126 ^ x20 ;
  assign n149 = x5 & ~n72 ;
  assign n150 = n107 & n149 ;
  assign n148 = x5 & ~n100 ;
  assign n151 = n150 ^ n148 ;
  assign n145 = x5 & n93 ;
  assign n146 = n145 ^ x5 ;
  assign n147 = n146 ^ x5 ;
  assign n152 = n151 ^ n147 ;
  assign n142 = x5 & n80 ;
  assign n143 = n142 ^ x5 ;
  assign n144 = n67 & n143 ;
  assign n153 = n152 ^ n144 ;
  assign n136 = x13 & ~n72 ;
  assign n137 = n107 & n136 ;
  assign n135 = x13 & ~n100 ;
  assign n138 = n137 ^ n135 ;
  assign n132 = x13 & n93 ;
  assign n133 = n132 ^ x13 ;
  assign n134 = n133 ^ x13 ;
  assign n139 = n138 ^ n134 ;
  assign n129 = x13 & n80 ;
  assign n130 = n129 ^ x13 ;
  assign n131 = n67 & n130 ;
  assign n140 = n139 ^ n131 ;
  assign n141 = n140 ^ x13 ;
  assign n154 = n153 ^ n141 ;
  assign n160 = n154 ^ x21 ;
  assign n161 = n128 & n160 ;
  assign n162 = n161 ^ n128 ;
  assign n163 = n162 ^ n160 ;
  assign n184 = x6 & ~n72 ;
  assign n185 = n107 & n184 ;
  assign n183 = x6 & ~n100 ;
  assign n186 = n185 ^ n183 ;
  assign n180 = x6 & n93 ;
  assign n181 = n180 ^ x6 ;
  assign n182 = n181 ^ x6 ;
  assign n187 = n186 ^ n182 ;
  assign n177 = x6 & n80 ;
  assign n178 = n177 ^ x6 ;
  assign n179 = n67 & n178 ;
  assign n188 = n187 ^ n179 ;
  assign n171 = x14 & ~n72 ;
  assign n172 = n107 & n171 ;
  assign n170 = x14 & ~n100 ;
  assign n173 = n172 ^ n170 ;
  assign n167 = x14 & n93 ;
  assign n168 = n167 ^ x14 ;
  assign n169 = n168 ^ x14 ;
  assign n174 = n173 ^ n169 ;
  assign n164 = x14 & n80 ;
  assign n165 = n164 ^ x14 ;
  assign n166 = n67 & n165 ;
  assign n175 = n174 ^ n166 ;
  assign n176 = n175 ^ x14 ;
  assign n189 = n188 ^ n176 ;
  assign n192 = n189 ^ x22 ;
  assign n212 = x7 & ~n72 ;
  assign n213 = n107 & n212 ;
  assign n211 = x7 & n100 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ x7 ;
  assign n208 = x7 & n93 ;
  assign n209 = n208 ^ x7 ;
  assign n210 = n209 ^ x7 ;
  assign n216 = n215 ^ n210 ;
  assign n205 = x7 & n80 ;
  assign n206 = n205 ^ x7 ;
  assign n207 = n67 & n206 ;
  assign n217 = n216 ^ n207 ;
  assign n200 = x15 & ~n72 ;
  assign n201 = n107 & n200 ;
  assign n199 = x15 & n100 ;
  assign n202 = n201 ^ n199 ;
  assign n196 = x15 & n93 ;
  assign n197 = n196 ^ x15 ;
  assign n198 = n197 ^ x15 ;
  assign n203 = n202 ^ n198 ;
  assign n193 = x15 & n80 ;
  assign n194 = n193 ^ x15 ;
  assign n195 = n67 & n194 ;
  assign n204 = n203 ^ n195 ;
  assign n218 = n217 ^ n204 ;
  assign n347 = n218 ^ x23 ;
  assign n348 = n192 & n347 ;
  assign n349 = n348 ^ n192 ;
  assign n350 = n349 ^ n347 ;
  assign n351 = n163 & n350 ;
  assign n352 = n351 ^ n163 ;
  assign n353 = n352 ^ n350 ;
  assign n354 = n343 & n353 ;
  assign n355 = n354 ^ n343 ;
  assign n356 = n355 ^ n353 ;
  assign n413 = x16 & n356 ;
  assign n414 = n413 ^ x16 ;
  assign n415 = n414 ^ x16 ;
  assign n420 = n419 ^ n415 ;
  assign n219 = x23 & n218 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = n192 & n220 ;
  assign n222 = n221 ^ n220 ;
  assign n190 = x22 & n189 ;
  assign n191 = n190 ^ n189 ;
  assign n223 = n222 ^ n191 ;
  assign n224 = n163 & n223 ;
  assign n225 = n224 ^ n223 ;
  assign n155 = x21 & n154 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n128 & n156 ;
  assign n158 = n157 ^ n156 ;
  assign n127 = ~x20 & n126 ;
  assign n159 = n158 ^ n127 ;
  assign n226 = n225 ^ n159 ;
  assign n410 = x16 & n343 ;
  assign n411 = n410 ^ x16 ;
  assign n412 = n226 & n411 ;
  assign n421 = n420 ^ n412 ;
  assign n721 = n421 ^ x16 ;
  assign n404 = n252 & ~n283 ;
  assign n405 = n370 & n404 ;
  assign n403 = n252 & ~n363 ;
  assign n406 = n405 ^ n403 ;
  assign n400 = n252 & n356 ;
  assign n401 = n400 ^ n252 ;
  assign n402 = n401 ^ n252 ;
  assign n407 = n406 ^ n402 ;
  assign n397 = n252 & n343 ;
  assign n398 = n397 ^ n252 ;
  assign n399 = n226 & n398 ;
  assign n408 = n407 ^ n399 ;
  assign n722 = n721 ^ n408 ;
  assign n724 = n722 ^ x24 ;
  assign n445 = x17 & ~n283 ;
  assign n446 = n370 & n445 ;
  assign n444 = x17 & ~n363 ;
  assign n447 = n446 ^ n444 ;
  assign n441 = x17 & n356 ;
  assign n442 = n441 ^ x17 ;
  assign n443 = n442 ^ x17 ;
  assign n448 = n447 ^ n443 ;
  assign n438 = x17 & n343 ;
  assign n439 = n438 ^ x17 ;
  assign n440 = n226 & n439 ;
  assign n449 = n448 ^ n440 ;
  assign n725 = n449 ^ x17 ;
  assign n432 = n279 & ~n283 ;
  assign n433 = n370 & n432 ;
  assign n431 = n279 & ~n363 ;
  assign n434 = n433 ^ n431 ;
  assign n428 = n279 & n356 ;
  assign n429 = n428 ^ n279 ;
  assign n430 = n429 ^ n279 ;
  assign n435 = n434 ^ n430 ;
  assign n425 = n279 & n343 ;
  assign n426 = n425 ^ n279 ;
  assign n427 = n226 & n426 ;
  assign n436 = n435 ^ n427 ;
  assign n726 = n725 ^ n436 ;
  assign n730 = n726 ^ x25 ;
  assign n731 = n724 & n730 ;
  assign n732 = n731 ^ n724 ;
  assign n733 = n732 ^ n730 ;
  assign n482 = x18 & ~n283 ;
  assign n483 = n370 & n482 ;
  assign n481 = x18 & ~n363 ;
  assign n484 = n483 ^ n481 ;
  assign n478 = x18 & n356 ;
  assign n479 = n478 ^ x18 ;
  assign n480 = n479 ^ x18 ;
  assign n485 = n484 ^ n480 ;
  assign n475 = x18 & n343 ;
  assign n476 = n475 ^ x18 ;
  assign n477 = n226 & n476 ;
  assign n486 = n485 ^ n477 ;
  assign n734 = n486 ^ x18 ;
  assign n469 = ~n283 & n309 ;
  assign n470 = n370 & n469 ;
  assign n468 = n309 & ~n363 ;
  assign n471 = n470 ^ n468 ;
  assign n465 = n309 & n356 ;
  assign n466 = n465 ^ n309 ;
  assign n467 = n466 ^ n309 ;
  assign n472 = n471 ^ n467 ;
  assign n462 = n309 & n343 ;
  assign n463 = n462 ^ n309 ;
  assign n464 = n226 & n463 ;
  assign n473 = n472 ^ n464 ;
  assign n735 = n734 ^ n473 ;
  assign n737 = n735 ^ x26 ;
  assign n512 = x19 & ~n283 ;
  assign n513 = n370 & n512 ;
  assign n511 = x19 & ~n363 ;
  assign n514 = n513 ^ n511 ;
  assign n508 = x19 & n356 ;
  assign n509 = n508 ^ x19 ;
  assign n510 = n509 ^ x19 ;
  assign n515 = n514 ^ n510 ;
  assign n505 = x19 & n343 ;
  assign n506 = n505 ^ x19 ;
  assign n507 = n226 & n506 ;
  assign n516 = n515 ^ n507 ;
  assign n738 = n516 ^ x19 ;
  assign n499 = ~n283 & n336 ;
  assign n500 = n370 & n499 ;
  assign n498 = n336 & ~n363 ;
  assign n501 = n500 ^ n498 ;
  assign n495 = n336 & n356 ;
  assign n496 = n495 ^ n336 ;
  assign n497 = n496 ^ n336 ;
  assign n502 = n501 ^ n497 ;
  assign n492 = n336 & n343 ;
  assign n493 = n492 ^ n336 ;
  assign n494 = n226 & n493 ;
  assign n503 = n502 ^ n494 ;
  assign n739 = n738 ^ n503 ;
  assign n748 = n739 ^ x27 ;
  assign n749 = n737 & n748 ;
  assign n750 = n749 ^ n737 ;
  assign n751 = n750 ^ n748 ;
  assign n752 = n733 & n751 ;
  assign n753 = n752 ^ n733 ;
  assign n754 = n753 ^ n751 ;
  assign n384 = x20 & ~n283 ;
  assign n385 = n370 & n384 ;
  assign n383 = x20 & ~n363 ;
  assign n386 = n385 ^ n383 ;
  assign n380 = x20 & n356 ;
  assign n381 = n380 ^ x20 ;
  assign n382 = n381 ^ x20 ;
  assign n387 = n386 ^ n382 ;
  assign n377 = x20 & n343 ;
  assign n378 = n377 ^ x20 ;
  assign n379 = n226 & n378 ;
  assign n388 = n387 ^ n379 ;
  assign n719 = n388 ^ x20 ;
  assign n371 = n126 & ~n283 ;
  assign n372 = n370 & n371 ;
  assign n364 = n126 & ~n363 ;
  assign n373 = n372 ^ n364 ;
  assign n357 = n126 & n356 ;
  assign n358 = n357 ^ n126 ;
  assign n359 = n358 ^ n126 ;
  assign n374 = n373 ^ n359 ;
  assign n344 = n126 & n343 ;
  assign n345 = n344 ^ n126 ;
  assign n346 = n226 & n345 ;
  assign n375 = n374 ^ n346 ;
  assign n720 = n719 ^ n375 ;
  assign n756 = n720 ^ x28 ;
  assign n559 = x21 & ~n283 ;
  assign n560 = n370 & n559 ;
  assign n558 = x21 & ~n363 ;
  assign n561 = n560 ^ n558 ;
  assign n555 = x21 & n356 ;
  assign n556 = n555 ^ x21 ;
  assign n557 = n556 ^ x21 ;
  assign n562 = n561 ^ n557 ;
  assign n552 = x21 & n343 ;
  assign n553 = n552 ^ x21 ;
  assign n554 = n226 & n553 ;
  assign n563 = n562 ^ n554 ;
  assign n757 = n563 ^ x21 ;
  assign n546 = n154 & ~n283 ;
  assign n547 = n370 & n546 ;
  assign n545 = n154 & ~n363 ;
  assign n548 = n547 ^ n545 ;
  assign n542 = n154 & n356 ;
  assign n543 = n542 ^ n154 ;
  assign n544 = n543 ^ n154 ;
  assign n549 = n548 ^ n544 ;
  assign n539 = n154 & n343 ;
  assign n540 = n539 ^ n154 ;
  assign n541 = n226 & n540 ;
  assign n550 = n549 ^ n541 ;
  assign n758 = n757 ^ n550 ;
  assign n764 = n758 ^ x29 ;
  assign n765 = n756 & n764 ;
  assign n766 = n765 ^ n756 ;
  assign n767 = n766 ^ n764 ;
  assign n649 = x22 & ~n283 ;
  assign n650 = n370 & n649 ;
  assign n648 = x22 & ~n363 ;
  assign n651 = n650 ^ n648 ;
  assign n645 = x22 & n356 ;
  assign n646 = n645 ^ x22 ;
  assign n647 = n646 ^ x22 ;
  assign n652 = n651 ^ n647 ;
  assign n642 = x22 & n343 ;
  assign n643 = n642 ^ x22 ;
  assign n644 = n226 & n643 ;
  assign n653 = n652 ^ n644 ;
  assign n805 = n653 ^ x22 ;
  assign n632 = n189 & ~n283 ;
  assign n633 = n370 & n632 ;
  assign n631 = n189 & ~n363 ;
  assign n634 = n633 ^ n631 ;
  assign n628 = n189 & n356 ;
  assign n629 = n628 ^ n189 ;
  assign n630 = n629 ^ n189 ;
  assign n635 = n634 ^ n630 ;
  assign n625 = n189 & n343 ;
  assign n626 = n625 ^ n189 ;
  assign n627 = n226 & n626 ;
  assign n636 = n635 ^ n627 ;
  assign n825 = n805 ^ n636 ;
  assign n826 = n825 ^ x30 ;
  assign n696 = x23 & ~n283 ;
  assign n697 = n370 & n696 ;
  assign n695 = x23 & ~n363 ;
  assign n698 = n697 ^ n695 ;
  assign n692 = x23 & n356 ;
  assign n693 = n692 ^ x23 ;
  assign n694 = n693 ^ x23 ;
  assign n699 = n698 ^ n694 ;
  assign n689 = x23 & n343 ;
  assign n690 = n689 ^ x23 ;
  assign n691 = n226 & n690 ;
  assign n700 = n699 ^ n691 ;
  assign n827 = n700 ^ x23 ;
  assign n683 = n218 & ~n283 ;
  assign n684 = n370 & n683 ;
  assign n682 = n218 & ~n363 ;
  assign n685 = n684 ^ n682 ;
  assign n679 = n218 & n356 ;
  assign n680 = n679 ^ n218 ;
  assign n681 = n680 ^ n218 ;
  assign n686 = n685 ^ n681 ;
  assign n676 = n218 & n343 ;
  assign n677 = n676 ^ n218 ;
  assign n678 = n226 & n677 ;
  assign n687 = n686 ^ n678 ;
  assign n828 = n827 ^ n687 ;
  assign n829 = n828 ^ x31 ;
  assign n830 = n826 & n829 ;
  assign n831 = n830 ^ n826 ;
  assign n832 = n831 ^ n829 ;
  assign n833 = n767 & n832 ;
  assign n834 = n833 ^ n767 ;
  assign n835 = n834 ^ n832 ;
  assign n836 = n754 & n835 ;
  assign n837 = n836 ^ n754 ;
  assign n838 = n837 ^ n835 ;
  assign n810 = x22 & ~x30 ;
  assign n814 = ~n356 & n810 ;
  assign n579 = ~n283 & n370 ;
  assign n580 = n579 ^ n363 ;
  assign n813 = ~n580 & n810 ;
  assign n815 = n814 ^ n813 ;
  assign n811 = ~n343 & n810 ;
  assign n812 = n226 & n811 ;
  assign n816 = n815 ^ n812 ;
  assign n788 = x23 & ~x31 ;
  assign n796 = ~n283 & n788 ;
  assign n797 = n370 & n796 ;
  assign n795 = ~n363 & n788 ;
  assign n798 = n797 ^ n795 ;
  assign n792 = n356 & n788 ;
  assign n793 = n792 ^ n788 ;
  assign n794 = n793 ^ n788 ;
  assign n799 = n798 ^ n794 ;
  assign n789 = n343 & n788 ;
  assign n790 = n789 ^ n788 ;
  assign n791 = n226 & n790 ;
  assign n800 = n799 ^ n791 ;
  assign n801 = n800 ^ n788 ;
  assign n775 = ~x31 & n218 ;
  assign n783 = ~n283 & n775 ;
  assign n784 = n370 & n783 ;
  assign n782 = ~n363 & n775 ;
  assign n785 = n784 ^ n782 ;
  assign n779 = n356 & n775 ;
  assign n780 = n779 ^ n775 ;
  assign n781 = n780 ^ n775 ;
  assign n786 = n785 ^ n781 ;
  assign n776 = n343 & n775 ;
  assign n777 = n776 ^ n775 ;
  assign n778 = n226 & n777 ;
  assign n787 = n786 ^ n778 ;
  assign n802 = n801 ^ n787 ;
  assign n807 = n636 & n802 ;
  assign n806 = n802 & n805 ;
  assign n808 = n807 ^ n806 ;
  assign n803 = x30 & n802 ;
  assign n804 = n803 ^ n802 ;
  assign n809 = n808 ^ n804 ;
  assign n817 = n816 ^ n809 ;
  assign n768 = ~x30 & n189 ;
  assign n772 = ~n580 & n768 ;
  assign n771 = n356 & n768 ;
  assign n773 = n772 ^ n771 ;
  assign n769 = ~n343 & n768 ;
  assign n770 = n226 & n769 ;
  assign n774 = n773 ^ n770 ;
  assign n818 = n817 ^ n774 ;
  assign n819 = n767 & n818 ;
  assign n820 = n819 ^ n818 ;
  assign n759 = x29 & n758 ;
  assign n760 = n759 ^ n758 ;
  assign n761 = n756 & n760 ;
  assign n762 = n761 ^ n760 ;
  assign n755 = ~x28 & n720 ;
  assign n763 = n762 ^ n755 ;
  assign n821 = n820 ^ n763 ;
  assign n822 = n754 & n821 ;
  assign n823 = n822 ^ n821 ;
  assign n740 = x27 & n739 ;
  assign n741 = n740 ^ n739 ;
  assign n742 = n737 & n741 ;
  assign n743 = n742 ^ n741 ;
  assign n736 = ~x26 & n735 ;
  assign n744 = n743 ^ n736 ;
  assign n745 = n733 & n744 ;
  assign n746 = n745 ^ n744 ;
  assign n727 = ~x25 & n726 ;
  assign n728 = ~n724 & n727 ;
  assign n723 = ~x24 & n722 ;
  assign n729 = n728 ^ n723 ;
  assign n747 = n746 ^ n729 ;
  assign n824 = n823 ^ n747 ;
  assign n839 = n838 ^ n824 ;
  assign n910 = x24 & n839 ;
  assign n911 = n910 ^ x24 ;
  assign n1340 = n911 ^ x24 ;
  assign n907 = n722 & n839 ;
  assign n908 = n907 ^ n722 ;
  assign n1341 = n1340 ^ n908 ;
  assign n1343 = n1341 ^ x32 ;
  assign n917 = x25 & n839 ;
  assign n918 = n917 ^ x25 ;
  assign n1344 = n918 ^ x25 ;
  assign n914 = n726 & n839 ;
  assign n915 = n914 ^ n726 ;
  assign n1345 = n1344 ^ n915 ;
  assign n1349 = n1345 ^ x33 ;
  assign n1350 = n1343 & n1349 ;
  assign n1351 = n1350 ^ n1343 ;
  assign n1352 = n1351 ^ n1349 ;
  assign n939 = x26 & n839 ;
  assign n940 = n939 ^ x26 ;
  assign n1353 = n940 ^ x26 ;
  assign n936 = n735 & n839 ;
  assign n937 = n936 ^ n735 ;
  assign n1354 = n1353 ^ n937 ;
  assign n1356 = n1354 ^ x34 ;
  assign n952 = x27 & n839 ;
  assign n953 = n952 ^ x27 ;
  assign n1362 = n953 ^ x27 ;
  assign n949 = n739 & n839 ;
  assign n950 = n949 ^ n739 ;
  assign n1363 = n1362 ^ n950 ;
  assign n1370 = n1363 ^ x35 ;
  assign n1371 = n1356 & n1370 ;
  assign n1372 = n1371 ^ n1356 ;
  assign n1373 = n1372 ^ n1370 ;
  assign n1374 = n1352 & n1373 ;
  assign n1375 = n1374 ^ n1352 ;
  assign n1376 = n1375 ^ n1373 ;
  assign n843 = x28 & n839 ;
  assign n844 = n843 ^ x28 ;
  assign n1338 = n844 ^ x28 ;
  assign n840 = n720 & n839 ;
  assign n841 = n840 ^ n720 ;
  assign n1339 = n1338 ^ n841 ;
  assign n1378 = n1339 ^ x36 ;
  assign n857 = x29 & n839 ;
  assign n858 = n857 ^ x29 ;
  assign n1384 = n858 ^ x29 ;
  assign n854 = n758 & n839 ;
  assign n855 = n854 ^ n758 ;
  assign n1385 = n1384 ^ n855 ;
  assign n1390 = n1385 ^ x37 ;
  assign n1391 = n1378 & n1390 ;
  assign n1392 = n1391 ^ n1378 ;
  assign n1393 = n1392 ^ n1390 ;
  assign n876 = x30 & n839 ;
  assign n877 = n876 ^ x30 ;
  assign n1424 = n877 ^ x30 ;
  assign n873 = n825 & n839 ;
  assign n874 = n873 ^ n825 ;
  assign n1425 = n1424 ^ n874 ;
  assign n1426 = n1425 ^ x38 ;
  assign n884 = x31 & n839 ;
  assign n885 = n884 ^ x31 ;
  assign n1427 = n885 ^ x31 ;
  assign n881 = n828 & n839 ;
  assign n882 = n881 ^ n828 ;
  assign n1428 = n1427 ^ n882 ;
  assign n1429 = n1428 ^ x39 ;
  assign n1430 = n1426 & n1429 ;
  assign n1431 = n1430 ^ n1426 ;
  assign n1432 = n1431 ^ n1429 ;
  assign n1433 = n1393 & n1432 ;
  assign n1434 = n1433 ^ n1393 ;
  assign n1435 = n1434 ^ n1432 ;
  assign n1436 = n1376 & n1435 ;
  assign n1437 = n1436 ^ n1376 ;
  assign n1438 = n1437 ^ n1435 ;
  assign n1414 = x30 & ~x38 ;
  assign n1415 = n839 & n1414 ;
  assign n1396 = ~x39 & n828 ;
  assign n1410 = n825 & n1396 ;
  assign n1411 = ~n839 & n1410 ;
  assign n1398 = x31 & ~x39 ;
  assign n1408 = x30 & n1398 ;
  assign n1409 = n839 & n1408 ;
  assign n1412 = n1411 ^ n1409 ;
  assign n1404 = x38 & n1396 ;
  assign n1405 = ~n839 & n1404 ;
  assign n1402 = x38 & n1398 ;
  assign n1403 = n839 & n1402 ;
  assign n1406 = n1405 ^ n1403 ;
  assign n1399 = ~n839 & n1398 ;
  assign n1400 = n1399 ^ n1398 ;
  assign n1397 = ~n839 & n1396 ;
  assign n1401 = n1400 ^ n1397 ;
  assign n1407 = n1406 ^ n1401 ;
  assign n1413 = n1412 ^ n1407 ;
  assign n1416 = n1415 ^ n1413 ;
  assign n1394 = ~x38 & n825 ;
  assign n1395 = ~n839 & n1394 ;
  assign n1417 = n1416 ^ n1395 ;
  assign n1418 = n1393 & n1417 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1381 = x29 & x37 ;
  assign n1382 = n839 & n1381 ;
  assign n1379 = x37 & n758 ;
  assign n1380 = ~n839 & n1379 ;
  assign n1383 = n1382 ^ n1380 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1387 = n1378 & n1386 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1377 = ~x36 & n1339 ;
  assign n1389 = n1388 ^ n1377 ;
  assign n1420 = n1419 ^ n1389 ;
  assign n1421 = n1376 & n1420 ;
  assign n1422 = n1421 ^ n1420 ;
  assign n1359 = x27 & x35 ;
  assign n1360 = n839 & n1359 ;
  assign n1357 = x35 & n739 ;
  assign n1358 = ~n839 & n1357 ;
  assign n1361 = n1360 ^ n1358 ;
  assign n1364 = n1363 ^ n1361 ;
  assign n1365 = n1356 & n1364 ;
  assign n1366 = n1365 ^ n1364 ;
  assign n1355 = ~x34 & n1354 ;
  assign n1367 = n1366 ^ n1355 ;
  assign n1368 = ~n1352 & n1367 ;
  assign n1346 = ~x33 & n1345 ;
  assign n1347 = ~n1343 & n1346 ;
  assign n1342 = ~x32 & n1341 ;
  assign n1348 = n1347 ^ n1342 ;
  assign n1369 = n1368 ^ n1348 ;
  assign n1423 = n1422 ^ n1369 ;
  assign n1439 = n1438 ^ n1423 ;
  assign n1497 = x32 & n1439 ;
  assign n1498 = n1497 ^ x32 ;
  assign n2198 = n1498 ^ x32 ;
  assign n1494 = n1341 & n1439 ;
  assign n1495 = n1494 ^ n1341 ;
  assign n2199 = n2198 ^ n1495 ;
  assign n2201 = n2199 ^ x40 ;
  assign n1506 = x33 & n1439 ;
  assign n1507 = n1506 ^ x33 ;
  assign n2202 = n1507 ^ x33 ;
  assign n1503 = n1345 & n1439 ;
  assign n1504 = n1503 ^ n1345 ;
  assign n2203 = n2202 ^ n1504 ;
  assign n2207 = n2203 ^ x41 ;
  assign n2208 = n2201 & n2207 ;
  assign n2209 = n2208 ^ n2201 ;
  assign n2210 = n2209 ^ n2207 ;
  assign n1516 = x34 & n1439 ;
  assign n1517 = n1516 ^ x34 ;
  assign n2211 = n1517 ^ x34 ;
  assign n1513 = n1354 & n1439 ;
  assign n1514 = n1513 ^ n1354 ;
  assign n2212 = n2211 ^ n1514 ;
  assign n2214 = n2212 ^ x42 ;
  assign n1527 = x35 & n1439 ;
  assign n1528 = n1527 ^ x35 ;
  assign n2220 = n1528 ^ x35 ;
  assign n1524 = n1363 & n1439 ;
  assign n1525 = n1524 ^ n1363 ;
  assign n2221 = n2220 ^ n1525 ;
  assign n2229 = n2221 ^ x43 ;
  assign n2230 = n2214 & n2229 ;
  assign n2231 = n2230 ^ n2214 ;
  assign n2232 = n2231 ^ n2229 ;
  assign n2233 = n2210 & n2232 ;
  assign n2234 = n2233 ^ n2210 ;
  assign n2235 = n2234 ^ n2232 ;
  assign n1443 = x36 & n1439 ;
  assign n1444 = n1443 ^ x36 ;
  assign n2196 = n1444 ^ x36 ;
  assign n1440 = n1339 & n1439 ;
  assign n1441 = n1440 ^ n1339 ;
  assign n2197 = n2196 ^ n1441 ;
  assign n2237 = n2197 ^ x44 ;
  assign n1453 = x37 & n1439 ;
  assign n1454 = n1453 ^ x37 ;
  assign n2243 = n1454 ^ x37 ;
  assign n1450 = n1385 & n1439 ;
  assign n1451 = n1450 ^ n1385 ;
  assign n2244 = n2243 ^ n1451 ;
  assign n2249 = n2244 ^ x45 ;
  assign n2250 = n2237 & n2249 ;
  assign n2251 = n2250 ^ n2237 ;
  assign n2252 = n2251 ^ n2249 ;
  assign n1470 = x38 & n1439 ;
  assign n1471 = n1470 ^ x38 ;
  assign n2283 = n1471 ^ x38 ;
  assign n1467 = n1425 & n1439 ;
  assign n1468 = n1467 ^ n1425 ;
  assign n2284 = n2283 ^ n1468 ;
  assign n2285 = n2284 ^ x46 ;
  assign n1479 = x39 & n1439 ;
  assign n1480 = n1479 ^ x39 ;
  assign n2286 = n1480 ^ x39 ;
  assign n1476 = n1428 & n1439 ;
  assign n1477 = n1476 ^ n1428 ;
  assign n2287 = n2286 ^ n1477 ;
  assign n2288 = n2287 ^ x47 ;
  assign n2289 = n2285 & n2288 ;
  assign n2290 = n2289 ^ n2285 ;
  assign n2291 = n2290 ^ n2288 ;
  assign n2292 = n2252 & n2291 ;
  assign n2293 = n2292 ^ n2252 ;
  assign n2294 = n2293 ^ n2291 ;
  assign n2295 = n2235 & n2294 ;
  assign n2296 = n2295 ^ n2235 ;
  assign n2297 = n2296 ^ n2294 ;
  assign n2273 = x38 & ~x46 ;
  assign n2274 = n1439 & n2273 ;
  assign n2255 = ~x47 & n1428 ;
  assign n2269 = n1425 & n2255 ;
  assign n2270 = ~n1439 & n2269 ;
  assign n2257 = x39 & ~x47 ;
  assign n2267 = x38 & n2257 ;
  assign n2268 = n1439 & n2267 ;
  assign n2271 = n2270 ^ n2268 ;
  assign n2263 = x46 & n2257 ;
  assign n2264 = n1439 & n2263 ;
  assign n2261 = x46 & n2255 ;
  assign n2262 = ~n1439 & n2261 ;
  assign n2265 = n2264 ^ n2262 ;
  assign n2258 = ~n1439 & n2257 ;
  assign n2259 = n2258 ^ n2257 ;
  assign n2256 = ~n1439 & n2255 ;
  assign n2260 = n2259 ^ n2256 ;
  assign n2266 = n2265 ^ n2260 ;
  assign n2272 = n2271 ^ n2266 ;
  assign n2275 = n2274 ^ n2272 ;
  assign n2253 = ~x46 & n1425 ;
  assign n2254 = ~n1439 & n2253 ;
  assign n2276 = n2275 ^ n2254 ;
  assign n2277 = n2252 & n2276 ;
  assign n2278 = n2277 ^ n2276 ;
  assign n2240 = x37 & x45 ;
  assign n2241 = n1439 & n2240 ;
  assign n2238 = x45 & n1385 ;
  assign n2239 = ~n1439 & n2238 ;
  assign n2242 = n2241 ^ n2239 ;
  assign n2245 = n2244 ^ n2242 ;
  assign n2246 = n2237 & n2245 ;
  assign n2247 = n2246 ^ n2245 ;
  assign n2236 = ~x44 & n2197 ;
  assign n2248 = n2247 ^ n2236 ;
  assign n2279 = n2278 ^ n2248 ;
  assign n2280 = n2235 & n2279 ;
  assign n2281 = n2280 ^ n2279 ;
  assign n2217 = x35 & x43 ;
  assign n2218 = n1439 & n2217 ;
  assign n2215 = x43 & n1363 ;
  assign n2216 = ~n1439 & n2215 ;
  assign n2219 = n2218 ^ n2216 ;
  assign n2222 = n2221 ^ n2219 ;
  assign n2223 = n2214 & n2222 ;
  assign n2224 = n2223 ^ n2222 ;
  assign n2213 = ~x42 & n2212 ;
  assign n2225 = n2224 ^ n2213 ;
  assign n2226 = n2210 & n2225 ;
  assign n2227 = n2226 ^ n2225 ;
  assign n2204 = ~x41 & n2203 ;
  assign n2205 = ~n2201 & n2204 ;
  assign n2200 = ~x40 & n2199 ;
  assign n2206 = n2205 ^ n2200 ;
  assign n2228 = n2227 ^ n2206 ;
  assign n2282 = n2281 ^ n2228 ;
  assign n2298 = n2297 ^ n2282 ;
  assign n2377 = x42 & n2298 ;
  assign n2378 = n2377 ^ x42 ;
  assign n2374 = n2212 & n2298 ;
  assign n2375 = n2374 ^ n2212 ;
  assign n2376 = n2375 ^ n2212 ;
  assign n2379 = n2378 ^ n2376 ;
  assign n938 = n937 ^ n735 ;
  assign n941 = n940 ^ n938 ;
  assign n391 = ~n72 & n107 ;
  assign n392 = n391 ^ n100 ;
  assign n390 = n67 & ~n80 ;
  assign n393 = n392 ^ n390 ;
  assign n394 = n393 ^ n93 ;
  assign n460 = x2 & n394 ;
  assign n461 = n460 ^ n295 ;
  assign n409 = n408 ^ n252 ;
  assign n422 = n421 ^ n409 ;
  assign n395 = x0 & n394 ;
  assign n396 = n395 ^ n238 ;
  assign n424 = n422 ^ n396 ;
  assign n451 = x1 & n394 ;
  assign n452 = n451 ^ n265 ;
  assign n437 = n436 ^ n279 ;
  assign n450 = n449 ^ n437 ;
  assign n456 = n452 ^ n450 ;
  assign n457 = n424 & n456 ;
  assign n458 = n457 ^ n424 ;
  assign n459 = n458 ^ n456 ;
  assign n474 = n473 ^ n309 ;
  assign n487 = n486 ^ n474 ;
  assign n489 = n487 ^ n461 ;
  assign n504 = n503 ^ n336 ;
  assign n517 = n516 ^ n504 ;
  assign n490 = x3 & n394 ;
  assign n491 = n490 ^ n322 ;
  assign n526 = n517 ^ n491 ;
  assign n527 = n489 & n526 ;
  assign n528 = n527 ^ n489 ;
  assign n529 = n528 ^ n526 ;
  assign n530 = n459 & n529 ;
  assign n531 = n530 ^ n459 ;
  assign n532 = n531 ^ n529 ;
  assign n533 = x4 & n394 ;
  assign n534 = n533 ^ n112 ;
  assign n376 = n375 ^ n126 ;
  assign n389 = n388 ^ n376 ;
  assign n536 = n534 ^ n389 ;
  assign n551 = n550 ^ n154 ;
  assign n564 = n563 ^ n551 ;
  assign n537 = x5 & n394 ;
  assign n538 = n537 ^ n140 ;
  assign n570 = n564 ^ n538 ;
  assign n571 = n536 & n570 ;
  assign n572 = n571 ^ n536 ;
  assign n573 = n572 ^ n570 ;
  assign n637 = n636 ^ n189 ;
  assign n674 = n653 ^ n637 ;
  assign n574 = x6 & n394 ;
  assign n575 = n574 ^ n175 ;
  assign n675 = n674 ^ n575 ;
  assign n688 = n687 ^ n218 ;
  assign n701 = n700 ^ n688 ;
  assign n588 = x15 & ~n392 ;
  assign n589 = n588 ^ n196 ;
  assign n590 = n589 ^ n195 ;
  assign n585 = x7 & ~n392 ;
  assign n586 = n585 ^ n209 ;
  assign n587 = n586 ^ n207 ;
  assign n591 = n590 ^ n587 ;
  assign n702 = n701 ^ n591 ;
  assign n703 = n675 & n702 ;
  assign n704 = n703 ^ n675 ;
  assign n705 = n704 ^ n702 ;
  assign n706 = n573 & n705 ;
  assign n707 = n706 ^ n573 ;
  assign n708 = n707 ^ n705 ;
  assign n709 = n532 & n708 ;
  assign n710 = n709 ^ n532 ;
  assign n711 = n710 ^ n708 ;
  assign n659 = ~x22 & n575 ;
  assign n663 = ~n580 & n659 ;
  assign n662 = n356 & n659 ;
  assign n664 = n663 ^ n662 ;
  assign n660 = ~n343 & n659 ;
  assign n661 = n226 & n660 ;
  assign n665 = n664 ^ n661 ;
  assign n606 = ~x23 & n591 ;
  assign n614 = ~n283 & n606 ;
  assign n615 = n370 & n614 ;
  assign n613 = ~n363 & n606 ;
  assign n616 = n615 ^ n613 ;
  assign n610 = n356 & n606 ;
  assign n611 = n610 ^ n606 ;
  assign n612 = n611 ^ n606 ;
  assign n617 = n616 ^ n612 ;
  assign n607 = n343 & n606 ;
  assign n608 = n607 ^ n606 ;
  assign n609 = n226 & n608 ;
  assign n618 = n617 ^ n609 ;
  assign n592 = ~n218 & n591 ;
  assign n600 = ~n283 & n592 ;
  assign n601 = n370 & n600 ;
  assign n599 = ~n363 & n592 ;
  assign n602 = n601 ^ n599 ;
  assign n596 = n356 & n592 ;
  assign n597 = n596 ^ n592 ;
  assign n598 = n597 ^ n592 ;
  assign n603 = n602 ^ n598 ;
  assign n593 = n343 & n592 ;
  assign n594 = n593 ^ n592 ;
  assign n595 = n226 & n594 ;
  assign n604 = n603 ^ n595 ;
  assign n605 = n604 ^ n592 ;
  assign n619 = n618 ^ n605 ;
  assign n621 = n226 & n343 ;
  assign n622 = n621 ^ n226 ;
  assign n623 = n622 ^ n580 ;
  assign n624 = n623 ^ n356 ;
  assign n654 = n653 ^ n624 ;
  assign n655 = n619 & n654 ;
  assign n656 = n655 ^ n619 ;
  assign n638 = n637 ^ n624 ;
  assign n639 = n619 & n638 ;
  assign n640 = n639 ^ n619 ;
  assign n641 = n640 ^ n619 ;
  assign n657 = n656 ^ n641 ;
  assign n620 = n575 & n619 ;
  assign n658 = n657 ^ n620 ;
  assign n666 = n665 ^ n658 ;
  assign n576 = ~n189 & n575 ;
  assign n582 = ~n356 & n576 ;
  assign n581 = n576 & ~n580 ;
  assign n583 = n582 ^ n581 ;
  assign n577 = ~n343 & n576 ;
  assign n578 = n226 & n577 ;
  assign n584 = n583 ^ n578 ;
  assign n667 = n666 ^ n584 ;
  assign n668 = n573 & n667 ;
  assign n669 = n668 ^ n667 ;
  assign n565 = n538 & n564 ;
  assign n566 = n565 ^ n538 ;
  assign n567 = n536 & n566 ;
  assign n568 = n567 ^ n566 ;
  assign n535 = ~n389 & n534 ;
  assign n569 = n568 ^ n535 ;
  assign n670 = n669 ^ n569 ;
  assign n671 = n532 & n670 ;
  assign n672 = n671 ^ n670 ;
  assign n518 = n491 & n517 ;
  assign n519 = n518 ^ n491 ;
  assign n520 = n489 & n519 ;
  assign n521 = n520 ^ n519 ;
  assign n488 = n461 & ~n487 ;
  assign n522 = n521 ^ n488 ;
  assign n523 = n459 & n522 ;
  assign n524 = n523 ^ n522 ;
  assign n453 = ~n450 & n452 ;
  assign n454 = ~n424 & n453 ;
  assign n423 = n396 & ~n422 ;
  assign n455 = n454 ^ n423 ;
  assign n525 = n524 ^ n455 ;
  assign n673 = n672 ^ n525 ;
  assign n712 = n711 ^ n673 ;
  assign n933 = n461 & n712 ;
  assign n934 = n933 ^ n461 ;
  assign n930 = n487 & n712 ;
  assign n931 = n930 ^ n487 ;
  assign n932 = n931 ^ n487 ;
  assign n935 = n934 ^ n932 ;
  assign n942 = n941 ^ n935 ;
  assign n946 = n491 & n712 ;
  assign n947 = n946 ^ n491 ;
  assign n943 = n517 & n712 ;
  assign n944 = n943 ^ n517 ;
  assign n945 = n944 ^ n517 ;
  assign n948 = n947 ^ n945 ;
  assign n951 = n950 ^ n739 ;
  assign n954 = n953 ^ n951 ;
  assign n984 = n948 & n954 ;
  assign n985 = n984 ^ n948 ;
  assign n986 = n942 & n985 ;
  assign n987 = n986 ^ n985 ;
  assign n983 = n935 & ~n941 ;
  assign n988 = n987 ^ n983 ;
  assign n909 = n908 ^ n722 ;
  assign n912 = n911 ^ n909 ;
  assign n904 = n396 & n712 ;
  assign n905 = n904 ^ n396 ;
  assign n901 = n422 & n712 ;
  assign n902 = n901 ^ n422 ;
  assign n903 = n902 ^ n422 ;
  assign n906 = n905 ^ n903 ;
  assign n913 = n912 ^ n906 ;
  assign n923 = n452 & n712 ;
  assign n924 = n923 ^ n452 ;
  assign n920 = n450 & n712 ;
  assign n921 = n920 ^ n450 ;
  assign n922 = n921 ^ n450 ;
  assign n925 = n924 ^ n922 ;
  assign n916 = n915 ^ n726 ;
  assign n919 = n918 ^ n916 ;
  assign n926 = n925 ^ n919 ;
  assign n927 = n913 & n926 ;
  assign n928 = n927 ^ n913 ;
  assign n929 = n928 ^ n926 ;
  assign n1071 = ~n929 & n941 ;
  assign n1072 = n988 & n1071 ;
  assign n979 = ~n919 & n925 ;
  assign n980 = ~n913 & n979 ;
  assign n978 = n906 & ~n912 ;
  assign n981 = n980 ^ n978 ;
  assign n1070 = n941 & n981 ;
  assign n1073 = n1072 ^ n1070 ;
  assign n1074 = n1073 ^ n941 ;
  assign n955 = n954 ^ n948 ;
  assign n956 = n942 & n955 ;
  assign n957 = n956 ^ n942 ;
  assign n958 = n957 ^ n955 ;
  assign n959 = n929 & n958 ;
  assign n960 = n959 ^ n929 ;
  assign n961 = n960 ^ n958 ;
  assign n842 = n841 ^ n720 ;
  assign n845 = n844 ^ n842 ;
  assign n716 = n534 & n712 ;
  assign n717 = n716 ^ n534 ;
  assign n713 = n389 & n712 ;
  assign n714 = n713 ^ n389 ;
  assign n715 = n714 ^ n389 ;
  assign n718 = n717 ^ n715 ;
  assign n847 = n845 ^ n718 ;
  assign n856 = n855 ^ n758 ;
  assign n859 = n858 ^ n856 ;
  assign n851 = n538 & n712 ;
  assign n852 = n851 ^ n538 ;
  assign n848 = n564 & n712 ;
  assign n849 = n848 ^ n564 ;
  assign n850 = n849 ^ n564 ;
  assign n853 = n852 ^ n850 ;
  assign n863 = n859 ^ n853 ;
  assign n864 = n847 & n863 ;
  assign n865 = n864 ^ n847 ;
  assign n866 = n865 ^ n863 ;
  assign n875 = n874 ^ n825 ;
  assign n878 = n877 ^ n875 ;
  assign n870 = n575 & n712 ;
  assign n871 = n870 ^ n575 ;
  assign n867 = n674 & n712 ;
  assign n868 = n867 ^ n674 ;
  assign n869 = n868 ^ n674 ;
  assign n872 = n871 ^ n869 ;
  assign n880 = n878 ^ n872 ;
  assign n890 = n591 & n712 ;
  assign n891 = n890 ^ n591 ;
  assign n887 = n701 & n712 ;
  assign n888 = n887 ^ n701 ;
  assign n889 = n888 ^ n701 ;
  assign n892 = n891 ^ n889 ;
  assign n883 = n882 ^ n828 ;
  assign n886 = n885 ^ n883 ;
  assign n965 = n892 ^ n886 ;
  assign n966 = n880 & n965 ;
  assign n967 = n966 ^ n880 ;
  assign n968 = n967 ^ n965 ;
  assign n969 = n866 & n968 ;
  assign n970 = n969 ^ n866 ;
  assign n971 = n970 ^ n968 ;
  assign n972 = n961 & n971 ;
  assign n973 = n972 ^ n961 ;
  assign n974 = n973 ^ n971 ;
  assign n1067 = n941 & n974 ;
  assign n1068 = n1067 ^ n941 ;
  assign n1069 = n1068 ^ n941 ;
  assign n1075 = n1074 ^ n1069 ;
  assign n893 = n886 & n892 ;
  assign n894 = n893 ^ n892 ;
  assign n895 = n880 & n894 ;
  assign n896 = n895 ^ n894 ;
  assign n879 = n872 & ~n878 ;
  assign n897 = n896 ^ n879 ;
  assign n898 = n866 & n897 ;
  assign n899 = n898 ^ n897 ;
  assign n860 = n853 & ~n859 ;
  assign n861 = ~n847 & n860 ;
  assign n846 = n718 & ~n845 ;
  assign n862 = n861 ^ n846 ;
  assign n900 = n899 ^ n862 ;
  assign n1064 = n941 & n961 ;
  assign n1065 = n1064 ^ n941 ;
  assign n1066 = n900 & n1065 ;
  assign n1076 = n1075 ^ n1066 ;
  assign n1519 = n1076 ^ n941 ;
  assign n1057 = ~n929 & n935 ;
  assign n1058 = n988 & n1057 ;
  assign n1056 = n935 & n981 ;
  assign n1059 = n1058 ^ n1056 ;
  assign n1060 = n1059 ^ n935 ;
  assign n1053 = n935 & n974 ;
  assign n1054 = n1053 ^ n935 ;
  assign n1055 = n1054 ^ n935 ;
  assign n1061 = n1060 ^ n1055 ;
  assign n1050 = n935 & n961 ;
  assign n1051 = n1050 ^ n935 ;
  assign n1052 = n900 & n1051 ;
  assign n1062 = n1061 ^ n1052 ;
  assign n1520 = n1519 ^ n1062 ;
  assign n1515 = n1514 ^ n1354 ;
  assign n1518 = n1517 ^ n1515 ;
  assign n1521 = n1520 ^ n1518 ;
  assign n1102 = ~n929 & n954 ;
  assign n1103 = n988 & n1102 ;
  assign n1101 = n954 & n981 ;
  assign n1104 = n1103 ^ n1101 ;
  assign n1105 = n1104 ^ n954 ;
  assign n1098 = n954 & n974 ;
  assign n1099 = n1098 ^ n954 ;
  assign n1100 = n1099 ^ n954 ;
  assign n1106 = n1105 ^ n1100 ;
  assign n1095 = n954 & n961 ;
  assign n1096 = n1095 ^ n954 ;
  assign n1097 = n900 & n1096 ;
  assign n1107 = n1106 ^ n1097 ;
  assign n1522 = n1107 ^ n954 ;
  assign n1088 = ~n929 & n948 ;
  assign n1089 = n988 & n1088 ;
  assign n1087 = n948 & n981 ;
  assign n1090 = n1089 ^ n1087 ;
  assign n1091 = n1090 ^ n948 ;
  assign n1084 = n948 & n974 ;
  assign n1085 = n1084 ^ n948 ;
  assign n1086 = n1085 ^ n948 ;
  assign n1092 = n1091 ^ n1086 ;
  assign n1081 = n948 & n961 ;
  assign n1082 = n1081 ^ n948 ;
  assign n1083 = n900 & n1082 ;
  assign n1093 = n1092 ^ n1083 ;
  assign n1523 = n1522 ^ n1093 ;
  assign n1526 = n1525 ^ n1363 ;
  assign n1529 = n1528 ^ n1526 ;
  assign n1558 = n1523 & n1529 ;
  assign n1559 = n1558 ^ n1523 ;
  assign n1560 = n1521 & n1559 ;
  assign n1561 = n1560 ^ n1559 ;
  assign n1557 = ~n1518 & n1520 ;
  assign n1562 = n1561 ^ n1557 ;
  assign n1496 = n1495 ^ n1341 ;
  assign n1499 = n1498 ^ n1496 ;
  assign n1003 = n912 & ~n929 ;
  assign n1004 = n988 & n1003 ;
  assign n1002 = n912 & n981 ;
  assign n1005 = n1004 ^ n1002 ;
  assign n1006 = n1005 ^ n912 ;
  assign n999 = n912 & n974 ;
  assign n1000 = n999 ^ n912 ;
  assign n1001 = n1000 ^ n912 ;
  assign n1007 = n1006 ^ n1001 ;
  assign n996 = n912 & n961 ;
  assign n997 = n996 ^ n912 ;
  assign n998 = n900 & n997 ;
  assign n1008 = n1007 ^ n998 ;
  assign n1492 = n1008 ^ n912 ;
  assign n989 = n906 & ~n929 ;
  assign n990 = n988 & n989 ;
  assign n982 = n906 & n981 ;
  assign n991 = n990 ^ n982 ;
  assign n992 = n991 ^ n906 ;
  assign n975 = n906 & n974 ;
  assign n976 = n975 ^ n906 ;
  assign n977 = n976 ^ n906 ;
  assign n993 = n992 ^ n977 ;
  assign n962 = n906 & n961 ;
  assign n963 = n962 ^ n906 ;
  assign n964 = n900 & n963 ;
  assign n994 = n993 ^ n964 ;
  assign n1493 = n1492 ^ n994 ;
  assign n1500 = n1499 ^ n1493 ;
  assign n1505 = n1504 ^ n1345 ;
  assign n1508 = n1507 ^ n1505 ;
  assign n1034 = n919 & ~n929 ;
  assign n1035 = n988 & n1034 ;
  assign n1033 = n919 & n981 ;
  assign n1036 = n1035 ^ n1033 ;
  assign n1037 = n1036 ^ n919 ;
  assign n1030 = n919 & n974 ;
  assign n1031 = n1030 ^ n919 ;
  assign n1032 = n1031 ^ n919 ;
  assign n1038 = n1037 ^ n1032 ;
  assign n1027 = n919 & n961 ;
  assign n1028 = n1027 ^ n919 ;
  assign n1029 = n900 & n1028 ;
  assign n1039 = n1038 ^ n1029 ;
  assign n1501 = n1039 ^ n919 ;
  assign n1020 = n925 & ~n929 ;
  assign n1021 = n988 & n1020 ;
  assign n1019 = n925 & n981 ;
  assign n1022 = n1021 ^ n1019 ;
  assign n1023 = n1022 ^ n925 ;
  assign n1016 = n925 & n974 ;
  assign n1017 = n1016 ^ n925 ;
  assign n1018 = n1017 ^ n925 ;
  assign n1024 = n1023 ^ n1018 ;
  assign n1013 = n925 & n961 ;
  assign n1014 = n1013 ^ n925 ;
  assign n1015 = n900 & n1014 ;
  assign n1025 = n1024 ^ n1015 ;
  assign n1502 = n1501 ^ n1025 ;
  assign n1509 = n1508 ^ n1502 ;
  assign n1510 = n1500 & n1509 ;
  assign n1511 = n1510 ^ n1500 ;
  assign n1512 = n1511 ^ n1509 ;
  assign n1632 = ~n1512 & n1518 ;
  assign n1633 = n1562 & n1632 ;
  assign n1553 = n1502 & ~n1508 ;
  assign n1554 = ~n1500 & n1553 ;
  assign n1552 = n1493 & ~n1499 ;
  assign n1555 = n1554 ^ n1552 ;
  assign n1631 = n1518 & n1555 ;
  assign n1634 = n1633 ^ n1631 ;
  assign n1530 = n1529 ^ n1523 ;
  assign n1531 = n1521 & n1530 ;
  assign n1532 = n1531 ^ n1521 ;
  assign n1533 = n1532 ^ n1530 ;
  assign n1534 = n1512 & n1533 ;
  assign n1535 = n1534 ^ n1512 ;
  assign n1536 = n1535 ^ n1533 ;
  assign n1442 = n1441 ^ n1339 ;
  assign n1445 = n1444 ^ n1442 ;
  assign n1146 = n845 & ~n929 ;
  assign n1147 = n988 & n1146 ;
  assign n1145 = n845 & n981 ;
  assign n1148 = n1147 ^ n1145 ;
  assign n1149 = n1148 ^ n845 ;
  assign n1142 = n845 & n974 ;
  assign n1143 = n1142 ^ n845 ;
  assign n1144 = n1143 ^ n845 ;
  assign n1150 = n1149 ^ n1144 ;
  assign n1139 = n845 & n961 ;
  assign n1140 = n1139 ^ n845 ;
  assign n1141 = n900 & n1140 ;
  assign n1151 = n1150 ^ n1141 ;
  assign n1336 = n1151 ^ n845 ;
  assign n1132 = n718 & ~n929 ;
  assign n1133 = n988 & n1132 ;
  assign n1131 = n718 & n981 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1135 = n1134 ^ n718 ;
  assign n1128 = n718 & n974 ;
  assign n1129 = n1128 ^ n718 ;
  assign n1130 = n1129 ^ n718 ;
  assign n1136 = n1135 ^ n1130 ;
  assign n1125 = n718 & n961 ;
  assign n1126 = n1125 ^ n718 ;
  assign n1127 = n900 & n1126 ;
  assign n1137 = n1136 ^ n1127 ;
  assign n1337 = n1336 ^ n1137 ;
  assign n1447 = n1445 ^ n1337 ;
  assign n1452 = n1451 ^ n1385 ;
  assign n1455 = n1454 ^ n1452 ;
  assign n1177 = n859 & ~n929 ;
  assign n1178 = n988 & n1177 ;
  assign n1176 = n859 & n981 ;
  assign n1179 = n1178 ^ n1176 ;
  assign n1180 = n1179 ^ n859 ;
  assign n1173 = n859 & n974 ;
  assign n1174 = n1173 ^ n859 ;
  assign n1175 = n1174 ^ n859 ;
  assign n1181 = n1180 ^ n1175 ;
  assign n1170 = n859 & n961 ;
  assign n1171 = n1170 ^ n859 ;
  assign n1172 = n900 & n1171 ;
  assign n1182 = n1181 ^ n1172 ;
  assign n1448 = n1182 ^ n859 ;
  assign n1163 = n853 & ~n929 ;
  assign n1164 = n988 & n1163 ;
  assign n1162 = n853 & n981 ;
  assign n1165 = n1164 ^ n1162 ;
  assign n1166 = n1165 ^ n853 ;
  assign n1159 = n853 & n974 ;
  assign n1160 = n1159 ^ n853 ;
  assign n1161 = n1160 ^ n853 ;
  assign n1167 = n1166 ^ n1161 ;
  assign n1156 = n853 & n961 ;
  assign n1157 = n1156 ^ n853 ;
  assign n1158 = n900 & n1157 ;
  assign n1168 = n1167 ^ n1158 ;
  assign n1449 = n1448 ^ n1168 ;
  assign n1461 = n1455 ^ n1449 ;
  assign n1462 = n1447 & n1461 ;
  assign n1463 = n1462 ^ n1447 ;
  assign n1464 = n1463 ^ n1461 ;
  assign n1469 = n1468 ^ n1425 ;
  assign n1472 = n1471 ^ n1469 ;
  assign n1262 = n878 & ~n929 ;
  assign n1263 = n988 & n1262 ;
  assign n1261 = n878 & n981 ;
  assign n1264 = n1263 ^ n1261 ;
  assign n1265 = n1264 ^ n878 ;
  assign n1258 = n878 & n974 ;
  assign n1259 = n1258 ^ n878 ;
  assign n1260 = n1259 ^ n878 ;
  assign n1266 = n1265 ^ n1260 ;
  assign n1255 = n878 & n961 ;
  assign n1256 = n1255 ^ n878 ;
  assign n1257 = n900 & n1256 ;
  assign n1267 = n1266 ^ n1257 ;
  assign n1465 = n1267 ^ n878 ;
  assign n1244 = n872 & ~n929 ;
  assign n1245 = n988 & n1244 ;
  assign n1243 = n872 & n981 ;
  assign n1246 = n1245 ^ n1243 ;
  assign n1247 = n1246 ^ n872 ;
  assign n1240 = n872 & n974 ;
  assign n1241 = n1240 ^ n872 ;
  assign n1242 = n1241 ^ n872 ;
  assign n1248 = n1247 ^ n1242 ;
  assign n1237 = n872 & n961 ;
  assign n1238 = n1237 ^ n872 ;
  assign n1239 = n900 & n1238 ;
  assign n1249 = n1248 ^ n1239 ;
  assign n1466 = n1465 ^ n1249 ;
  assign n1475 = n1472 ^ n1466 ;
  assign n1312 = n886 & ~n929 ;
  assign n1313 = n988 & n1312 ;
  assign n1311 = n886 & n981 ;
  assign n1314 = n1313 ^ n1311 ;
  assign n1315 = n1314 ^ n886 ;
  assign n1308 = n886 & n974 ;
  assign n1309 = n1308 ^ n886 ;
  assign n1310 = n1309 ^ n886 ;
  assign n1316 = n1315 ^ n1310 ;
  assign n1305 = n886 & n961 ;
  assign n1306 = n1305 ^ n886 ;
  assign n1307 = n900 & n1306 ;
  assign n1317 = n1316 ^ n1307 ;
  assign n1482 = n1317 ^ n886 ;
  assign n1300 = n892 & n961 ;
  assign n1301 = n1300 ^ n892 ;
  assign n1302 = n900 & n1301 ;
  assign n1296 = n892 & n974 ;
  assign n1297 = n1296 ^ n892 ;
  assign n1298 = n1297 ^ n892 ;
  assign n1292 = n892 & ~n929 ;
  assign n1293 = n988 & n1292 ;
  assign n1291 = n892 & n981 ;
  assign n1294 = n1293 ^ n1291 ;
  assign n1295 = n1294 ^ n892 ;
  assign n1299 = n1298 ^ n1295 ;
  assign n1303 = n1302 ^ n1299 ;
  assign n1483 = n1482 ^ n1303 ;
  assign n1478 = n1477 ^ n1428 ;
  assign n1481 = n1480 ^ n1478 ;
  assign n1540 = n1483 ^ n1481 ;
  assign n1541 = n1475 & n1540 ;
  assign n1542 = n1541 ^ n1475 ;
  assign n1543 = n1542 ^ n1540 ;
  assign n1544 = n1464 & n1543 ;
  assign n1545 = n1544 ^ n1464 ;
  assign n1546 = n1545 ^ n1543 ;
  assign n1547 = n1536 & n1546 ;
  assign n1548 = n1547 ^ n1536 ;
  assign n1549 = n1548 ^ n1546 ;
  assign n1629 = n1518 & n1549 ;
  assign n1630 = n1629 ^ n1518 ;
  assign n1635 = n1634 ^ n1630 ;
  assign n1484 = n1481 & n1483 ;
  assign n1485 = n1484 ^ n1483 ;
  assign n1486 = n1475 & n1485 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1473 = n1466 & n1472 ;
  assign n1474 = n1473 ^ n1466 ;
  assign n1488 = n1487 ^ n1474 ;
  assign n1489 = n1464 & n1488 ;
  assign n1490 = n1489 ^ n1488 ;
  assign n1456 = n1449 & n1455 ;
  assign n1457 = n1456 ^ n1449 ;
  assign n1458 = n1447 & n1457 ;
  assign n1459 = n1458 ^ n1457 ;
  assign n1446 = n1337 & ~n1445 ;
  assign n1460 = n1459 ^ n1446 ;
  assign n1491 = n1490 ^ n1460 ;
  assign n1626 = n1518 & n1536 ;
  assign n1627 = n1626 ^ n1518 ;
  assign n1628 = n1491 & n1627 ;
  assign n1636 = n1635 ^ n1628 ;
  assign n2372 = n1636 ^ n1518 ;
  assign n1620 = ~n1512 & n1520 ;
  assign n1621 = n1562 & n1620 ;
  assign n1619 = n1520 & n1555 ;
  assign n1622 = n1621 ^ n1619 ;
  assign n1617 = n1520 & n1549 ;
  assign n1618 = n1617 ^ n1520 ;
  assign n1623 = n1622 ^ n1618 ;
  assign n1614 = n1520 & n1536 ;
  assign n1615 = n1614 ^ n1520 ;
  assign n1616 = n1491 & n1615 ;
  assign n1624 = n1623 ^ n1616 ;
  assign n2373 = n2372 ^ n1624 ;
  assign n2380 = n2379 ^ n2373 ;
  assign n1661 = ~n1512 & n1529 ;
  assign n1662 = n1562 & n1661 ;
  assign n1660 = n1529 & n1555 ;
  assign n1663 = n1662 ^ n1660 ;
  assign n1658 = n1529 & n1549 ;
  assign n1659 = n1658 ^ n1529 ;
  assign n1664 = n1663 ^ n1659 ;
  assign n1655 = n1529 & n1536 ;
  assign n1656 = n1655 ^ n1529 ;
  assign n1657 = n1491 & n1656 ;
  assign n1665 = n1664 ^ n1657 ;
  assign n2381 = n1665 ^ n1529 ;
  assign n1649 = ~n1512 & n1523 ;
  assign n1650 = n1562 & n1649 ;
  assign n1648 = n1523 & n1555 ;
  assign n1651 = n1650 ^ n1648 ;
  assign n1646 = n1523 & n1549 ;
  assign n1647 = n1646 ^ n1523 ;
  assign n1652 = n1651 ^ n1647 ;
  assign n1643 = n1523 & n1536 ;
  assign n1644 = n1643 ^ n1523 ;
  assign n1645 = n1491 & n1644 ;
  assign n1653 = n1652 ^ n1645 ;
  assign n2382 = n2381 ^ n1653 ;
  assign n2386 = x43 & n2298 ;
  assign n2387 = n2386 ^ x43 ;
  assign n2383 = n2221 & n2298 ;
  assign n2384 = n2383 ^ n2221 ;
  assign n2385 = n2384 ^ n2221 ;
  assign n2388 = n2387 ^ n2385 ;
  assign n2418 = n2382 & n2388 ;
  assign n2419 = n2418 ^ n2382 ;
  assign n2420 = n2380 & n2419 ;
  assign n2421 = n2420 ^ n2419 ;
  assign n2417 = n2373 & ~n2379 ;
  assign n2422 = n2421 ^ n2417 ;
  assign n2356 = x40 & n2298 ;
  assign n2357 = n2356 ^ x40 ;
  assign n2353 = n2199 & n2298 ;
  assign n2354 = n2353 ^ n2199 ;
  assign n2355 = n2354 ^ n2199 ;
  assign n2358 = n2357 ^ n2355 ;
  assign n1575 = n1499 & ~n1512 ;
  assign n1576 = n1562 & n1575 ;
  assign n1574 = n1499 & n1555 ;
  assign n1577 = n1576 ^ n1574 ;
  assign n1572 = n1499 & n1549 ;
  assign n1573 = n1572 ^ n1499 ;
  assign n1578 = n1577 ^ n1573 ;
  assign n1569 = n1499 & n1536 ;
  assign n1570 = n1569 ^ n1499 ;
  assign n1571 = n1491 & n1570 ;
  assign n1579 = n1578 ^ n1571 ;
  assign n2351 = n1579 ^ n1499 ;
  assign n1563 = n1493 & ~n1512 ;
  assign n1564 = n1562 & n1563 ;
  assign n1556 = n1493 & n1555 ;
  assign n1565 = n1564 ^ n1556 ;
  assign n1550 = n1493 & n1549 ;
  assign n1551 = n1550 ^ n1493 ;
  assign n1566 = n1565 ^ n1551 ;
  assign n1537 = n1493 & n1536 ;
  assign n1538 = n1537 ^ n1493 ;
  assign n1539 = n1491 & n1538 ;
  assign n1567 = n1566 ^ n1539 ;
  assign n2352 = n2351 ^ n1567 ;
  assign n2359 = n2358 ^ n2352 ;
  assign n2365 = x41 & n2298 ;
  assign n2366 = n2365 ^ x41 ;
  assign n2362 = n2203 & n2298 ;
  assign n2363 = n2362 ^ n2203 ;
  assign n2364 = n2363 ^ n2203 ;
  assign n2367 = n2366 ^ n2364 ;
  assign n1604 = n1508 & ~n1512 ;
  assign n1605 = n1562 & n1604 ;
  assign n1603 = n1508 & n1555 ;
  assign n1606 = n1605 ^ n1603 ;
  assign n1601 = n1508 & n1549 ;
  assign n1602 = n1601 ^ n1508 ;
  assign n1607 = n1606 ^ n1602 ;
  assign n1598 = n1508 & n1536 ;
  assign n1599 = n1598 ^ n1508 ;
  assign n1600 = n1491 & n1599 ;
  assign n1608 = n1607 ^ n1600 ;
  assign n2360 = n1608 ^ n1508 ;
  assign n1592 = n1502 & ~n1512 ;
  assign n1593 = n1562 & n1592 ;
  assign n1591 = n1502 & n1555 ;
  assign n1594 = n1593 ^ n1591 ;
  assign n1589 = n1502 & n1549 ;
  assign n1590 = n1589 ^ n1502 ;
  assign n1595 = n1594 ^ n1590 ;
  assign n1586 = n1502 & n1536 ;
  assign n1587 = n1586 ^ n1502 ;
  assign n1588 = n1491 & n1587 ;
  assign n1596 = n1595 ^ n1588 ;
  assign n2361 = n2360 ^ n1596 ;
  assign n2368 = n2367 ^ n2361 ;
  assign n2369 = n2359 & n2368 ;
  assign n2370 = n2369 ^ n2359 ;
  assign n2371 = n2370 ^ n2368 ;
  assign n2582 = n2358 & ~n2371 ;
  assign n2583 = n2422 & n2582 ;
  assign n2413 = n2361 & ~n2367 ;
  assign n2414 = ~n2359 & n2413 ;
  assign n2412 = n2352 & ~n2358 ;
  assign n2415 = n2414 ^ n2412 ;
  assign n2581 = n2358 & n2415 ;
  assign n2584 = n2583 ^ n2581 ;
  assign n2585 = n2584 ^ n2358 ;
  assign n2389 = n2388 ^ n2382 ;
  assign n2390 = n2380 & n2389 ;
  assign n2391 = n2390 ^ n2380 ;
  assign n2392 = n2391 ^ n2389 ;
  assign n2393 = n2371 & n2392 ;
  assign n2394 = n2393 ^ n2371 ;
  assign n2395 = n2394 ^ n2392 ;
  assign n2302 = x44 & n2298 ;
  assign n2303 = n2302 ^ x44 ;
  assign n2299 = n2197 & n2298 ;
  assign n2300 = n2299 ^ n2197 ;
  assign n2301 = n2300 ^ n2197 ;
  assign n2304 = n2303 ^ n2301 ;
  assign n1700 = n1445 & ~n1512 ;
  assign n1701 = n1562 & n1700 ;
  assign n1699 = n1445 & n1555 ;
  assign n1702 = n1701 ^ n1699 ;
  assign n1697 = n1445 & n1549 ;
  assign n1698 = n1697 ^ n1445 ;
  assign n1703 = n1702 ^ n1698 ;
  assign n1694 = n1445 & n1536 ;
  assign n1695 = n1694 ^ n1445 ;
  assign n1696 = n1491 & n1695 ;
  assign n1704 = n1703 ^ n1696 ;
  assign n2194 = n1704 ^ n1445 ;
  assign n1688 = n1337 & ~n1512 ;
  assign n1689 = n1562 & n1688 ;
  assign n1687 = n1337 & n1555 ;
  assign n1690 = n1689 ^ n1687 ;
  assign n1685 = n1337 & n1549 ;
  assign n1686 = n1685 ^ n1337 ;
  assign n1691 = n1690 ^ n1686 ;
  assign n1682 = n1337 & n1536 ;
  assign n1683 = n1682 ^ n1337 ;
  assign n1684 = n1491 & n1683 ;
  assign n1692 = n1691 ^ n1684 ;
  assign n2195 = n2194 ^ n1692 ;
  assign n2306 = n2304 ^ n2195 ;
  assign n2312 = x45 & n2298 ;
  assign n2313 = n2312 ^ x45 ;
  assign n2309 = n2244 & n2298 ;
  assign n2310 = n2309 ^ n2244 ;
  assign n2311 = n2310 ^ n2244 ;
  assign n2314 = n2313 ^ n2311 ;
  assign n1729 = n1455 & ~n1512 ;
  assign n1730 = n1562 & n1729 ;
  assign n1728 = n1455 & n1555 ;
  assign n1731 = n1730 ^ n1728 ;
  assign n1726 = n1455 & n1549 ;
  assign n1727 = n1726 ^ n1455 ;
  assign n1732 = n1731 ^ n1727 ;
  assign n1723 = n1455 & n1536 ;
  assign n1724 = n1723 ^ n1455 ;
  assign n1725 = n1491 & n1724 ;
  assign n1733 = n1732 ^ n1725 ;
  assign n2307 = n1733 ^ n1455 ;
  assign n1717 = n1449 & ~n1512 ;
  assign n1718 = n1562 & n1717 ;
  assign n1716 = n1449 & n1555 ;
  assign n1719 = n1718 ^ n1716 ;
  assign n1714 = n1449 & n1549 ;
  assign n1715 = n1714 ^ n1449 ;
  assign n1720 = n1719 ^ n1715 ;
  assign n1711 = n1449 & n1536 ;
  assign n1712 = n1711 ^ n1449 ;
  assign n1713 = n1491 & n1712 ;
  assign n1721 = n1720 ^ n1713 ;
  assign n2308 = n2307 ^ n1721 ;
  assign n2320 = n2314 ^ n2308 ;
  assign n2321 = n2306 & n2320 ;
  assign n2322 = n2321 ^ n2306 ;
  assign n2323 = n2322 ^ n2320 ;
  assign n2329 = x46 & n2298 ;
  assign n2330 = n2329 ^ x46 ;
  assign n2326 = n2284 & n2298 ;
  assign n2327 = n2326 ^ n2284 ;
  assign n2328 = n2327 ^ n2284 ;
  assign n2331 = n2330 ^ n2328 ;
  assign n1761 = n1472 & ~n1512 ;
  assign n1762 = n1562 & n1761 ;
  assign n1760 = n1472 & n1555 ;
  assign n1763 = n1762 ^ n1760 ;
  assign n1758 = n1472 & n1549 ;
  assign n1759 = n1758 ^ n1472 ;
  assign n1764 = n1763 ^ n1759 ;
  assign n1755 = n1472 & n1536 ;
  assign n1756 = n1755 ^ n1472 ;
  assign n1757 = n1491 & n1756 ;
  assign n1765 = n1764 ^ n1757 ;
  assign n2324 = n1765 ^ n1472 ;
  assign n1749 = n1466 & ~n1512 ;
  assign n1750 = n1562 & n1749 ;
  assign n1748 = n1466 & n1555 ;
  assign n1751 = n1750 ^ n1748 ;
  assign n1746 = n1466 & n1549 ;
  assign n1747 = n1746 ^ n1466 ;
  assign n1752 = n1751 ^ n1747 ;
  assign n1743 = n1466 & n1536 ;
  assign n1744 = n1743 ^ n1466 ;
  assign n1745 = n1491 & n1744 ;
  assign n1753 = n1752 ^ n1745 ;
  assign n2325 = n2324 ^ n1753 ;
  assign n2334 = n2331 ^ n2325 ;
  assign n2340 = x47 & n2298 ;
  assign n2341 = n2340 ^ x47 ;
  assign n2337 = n2287 & n2298 ;
  assign n2338 = n2337 ^ n2287 ;
  assign n2339 = n2338 ^ n2287 ;
  assign n2342 = n2341 ^ n2339 ;
  assign n1789 = n1481 & ~n1512 ;
  assign n1790 = n1562 & n1789 ;
  assign n1788 = n1481 & n1555 ;
  assign n1791 = n1790 ^ n1788 ;
  assign n1792 = n1791 ^ n1481 ;
  assign n1785 = n1481 & n1549 ;
  assign n1786 = n1785 ^ n1481 ;
  assign n1787 = n1786 ^ n1481 ;
  assign n1793 = n1792 ^ n1787 ;
  assign n1782 = n1481 & n1536 ;
  assign n1783 = n1782 ^ n1481 ;
  assign n1784 = n1491 & n1783 ;
  assign n1794 = n1793 ^ n1784 ;
  assign n2335 = n1794 ^ n1481 ;
  assign n1775 = n1483 & ~n1512 ;
  assign n1776 = n1562 & n1775 ;
  assign n1774 = n1483 & n1555 ;
  assign n1777 = n1776 ^ n1774 ;
  assign n1778 = n1777 ^ n1483 ;
  assign n1771 = n1483 & n1549 ;
  assign n1772 = n1771 ^ n1483 ;
  assign n1773 = n1772 ^ n1483 ;
  assign n1779 = n1778 ^ n1773 ;
  assign n1768 = n1483 & n1536 ;
  assign n1769 = n1768 ^ n1483 ;
  assign n1770 = n1491 & n1769 ;
  assign n1780 = n1779 ^ n1770 ;
  assign n2336 = n2335 ^ n1780 ;
  assign n2399 = n2342 ^ n2336 ;
  assign n2400 = n2334 & n2399 ;
  assign n2401 = n2400 ^ n2334 ;
  assign n2402 = n2401 ^ n2399 ;
  assign n2403 = n2323 & n2402 ;
  assign n2404 = n2403 ^ n2323 ;
  assign n2405 = n2404 ^ n2402 ;
  assign n2406 = n2395 & n2405 ;
  assign n2407 = n2406 ^ n2395 ;
  assign n2408 = n2407 ^ n2405 ;
  assign n2578 = n2358 & n2408 ;
  assign n2579 = n2578 ^ n2358 ;
  assign n2580 = n2579 ^ n2358 ;
  assign n2586 = n2585 ^ n2580 ;
  assign n2343 = n2336 & n2342 ;
  assign n2344 = n2343 ^ n2336 ;
  assign n2345 = n2334 & n2344 ;
  assign n2346 = n2345 ^ n2344 ;
  assign n2332 = n2325 & n2331 ;
  assign n2333 = n2332 ^ n2325 ;
  assign n2347 = n2346 ^ n2333 ;
  assign n2348 = n2323 & n2347 ;
  assign n2349 = n2348 ^ n2347 ;
  assign n2315 = n2308 & n2314 ;
  assign n2316 = n2315 ^ n2308 ;
  assign n2317 = n2306 & n2316 ;
  assign n2318 = n2317 ^ n2316 ;
  assign n2305 = n2195 & ~n2304 ;
  assign n2319 = n2318 ^ n2305 ;
  assign n2350 = n2349 ^ n2319 ;
  assign n2575 = n2358 & n2395 ;
  assign n2576 = n2575 ^ n2358 ;
  assign n2577 = n2350 & n2576 ;
  assign n2587 = n2586 ^ n2577 ;
  assign n2570 = n2352 & ~n2371 ;
  assign n2571 = n2422 & n2570 ;
  assign n2569 = n2352 & n2415 ;
  assign n2572 = n2571 ^ n2569 ;
  assign n2566 = n2352 & n2408 ;
  assign n2567 = n2566 ^ n2352 ;
  assign n2568 = n2567 ^ n2352 ;
  assign n2573 = n2572 ^ n2568 ;
  assign n2563 = n2352 & n2395 ;
  assign n2564 = n2563 ^ n2352 ;
  assign n2565 = n2350 & n2564 ;
  assign n2574 = n2573 ^ n2565 ;
  assign n2588 = n2587 ^ n2574 ;
  assign n1010 = n904 ^ n902 ;
  assign n995 = n994 ^ n906 ;
  assign n1009 = n1008 ^ n995 ;
  assign n1012 = n1010 ^ n1009 ;
  assign n1041 = n923 ^ n921 ;
  assign n1026 = n1025 ^ n925 ;
  assign n1040 = n1039 ^ n1026 ;
  assign n1045 = n1041 ^ n1040 ;
  assign n1046 = n1012 & n1045 ;
  assign n1047 = n1046 ^ n1012 ;
  assign n1048 = n1047 ^ n1045 ;
  assign n1063 = n1062 ^ n935 ;
  assign n1077 = n1076 ^ n1063 ;
  assign n1049 = n933 ^ n931 ;
  assign n1079 = n1077 ^ n1049 ;
  assign n1094 = n1093 ^ n948 ;
  assign n1108 = n1107 ^ n1094 ;
  assign n1080 = n946 ^ n944 ;
  assign n1117 = n1108 ^ n1080 ;
  assign n1118 = n1079 & n1117 ;
  assign n1119 = n1118 ^ n1079 ;
  assign n1120 = n1119 ^ n1117 ;
  assign n1121 = n1048 & n1120 ;
  assign n1122 = n1121 ^ n1048 ;
  assign n1123 = n1122 ^ n1120 ;
  assign n1138 = n1137 ^ n718 ;
  assign n1152 = n1151 ^ n1138 ;
  assign n1124 = n716 ^ n714 ;
  assign n1154 = n1152 ^ n1124 ;
  assign n1169 = n1168 ^ n853 ;
  assign n1183 = n1182 ^ n1169 ;
  assign n1155 = n851 ^ n849 ;
  assign n1189 = n1183 ^ n1155 ;
  assign n1190 = n1154 & n1189 ;
  assign n1191 = n1190 ^ n1154 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n1250 = n1249 ^ n872 ;
  assign n1289 = n1267 ^ n1250 ;
  assign n1200 = n870 ^ n868 ;
  assign n1290 = n1289 ^ n1200 ;
  assign n1304 = n1303 ^ n892 ;
  assign n1318 = n1317 ^ n1304 ;
  assign n1205 = n890 ^ n888 ;
  assign n1319 = n1318 ^ n1205 ;
  assign n1320 = n1290 & n1319 ;
  assign n1321 = n1320 ^ n1290 ;
  assign n1322 = n1321 ^ n1319 ;
  assign n1323 = n1192 & n1322 ;
  assign n1324 = n1323 ^ n1192 ;
  assign n1325 = n1324 ^ n1322 ;
  assign n1326 = n1123 & n1325 ;
  assign n1327 = n1326 ^ n1123 ;
  assign n1328 = n1327 ^ n1325 ;
  assign n1273 = ~n878 & n1200 ;
  assign n1277 = ~n961 & n1273 ;
  assign n1278 = n900 & n1277 ;
  assign n1275 = ~n971 & n1273 ;
  assign n1276 = ~n961 & n1275 ;
  assign n1279 = n1278 ^ n1276 ;
  assign n1195 = n929 & n988 ;
  assign n1196 = n1195 ^ n988 ;
  assign n1197 = n1196 ^ n981 ;
  assign n1274 = n1197 & n1273 ;
  assign n1280 = n1279 ^ n1274 ;
  assign n1220 = ~n892 & n1205 ;
  assign n1228 = ~n929 & n1220 ;
  assign n1229 = n988 & n1228 ;
  assign n1227 = n981 & n1220 ;
  assign n1230 = n1229 ^ n1227 ;
  assign n1231 = n1230 ^ n1220 ;
  assign n1224 = n974 & n1220 ;
  assign n1225 = n1224 ^ n1220 ;
  assign n1226 = n1225 ^ n1220 ;
  assign n1232 = n1231 ^ n1226 ;
  assign n1221 = n961 & n1220 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1223 = n900 & n1222 ;
  assign n1233 = n1232 ^ n1223 ;
  assign n1234 = n1233 ^ n1220 ;
  assign n1206 = ~n886 & n1205 ;
  assign n1214 = ~n929 & n1206 ;
  assign n1215 = n988 & n1214 ;
  assign n1213 = n981 & n1206 ;
  assign n1216 = n1215 ^ n1213 ;
  assign n1217 = n1216 ^ n1206 ;
  assign n1210 = n974 & n1206 ;
  assign n1211 = n1210 ^ n1206 ;
  assign n1212 = n1211 ^ n1206 ;
  assign n1218 = n1217 ^ n1212 ;
  assign n1207 = n961 & n1206 ;
  assign n1208 = n1207 ^ n1206 ;
  assign n1209 = n900 & n1208 ;
  assign n1219 = n1218 ^ n1209 ;
  assign n1235 = n1234 ^ n1219 ;
  assign n1193 = n900 & n961 ;
  assign n1194 = n1193 ^ n900 ;
  assign n1198 = n1197 ^ n1194 ;
  assign n1199 = n1198 ^ n974 ;
  assign n1268 = n1267 ^ n1199 ;
  assign n1269 = n1235 & n1268 ;
  assign n1270 = n1269 ^ n1235 ;
  assign n1251 = n1250 ^ n1199 ;
  assign n1252 = n1235 & n1251 ;
  assign n1253 = n1252 ^ n1235 ;
  assign n1254 = n1253 ^ n1235 ;
  assign n1271 = n1270 ^ n1254 ;
  assign n1236 = n1200 & n1235 ;
  assign n1272 = n1271 ^ n1236 ;
  assign n1281 = n1280 ^ n1272 ;
  assign n1201 = ~n872 & n1200 ;
  assign n1202 = n1199 & n1201 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1204 = n1203 ^ n1201 ;
  assign n1282 = n1281 ^ n1204 ;
  assign n1283 = n1192 & n1282 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1184 = n1155 & n1183 ;
  assign n1185 = n1184 ^ n1155 ;
  assign n1186 = n1154 & n1185 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1153 = n1124 & ~n1152 ;
  assign n1188 = n1187 ^ n1153 ;
  assign n1285 = n1284 ^ n1188 ;
  assign n1286 = n1123 & n1285 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1109 = n1080 & n1108 ;
  assign n1110 = n1109 ^ n1080 ;
  assign n1111 = n1079 & n1110 ;
  assign n1112 = n1111 ^ n1110 ;
  assign n1078 = n1049 & ~n1077 ;
  assign n1113 = n1112 ^ n1078 ;
  assign n1114 = n1048 & n1113 ;
  assign n1115 = n1114 ^ n1113 ;
  assign n1042 = ~n1040 & n1041 ;
  assign n1043 = ~n1012 & n1042 ;
  assign n1011 = ~n1009 & n1010 ;
  assign n1044 = n1043 ^ n1011 ;
  assign n1116 = n1115 ^ n1044 ;
  assign n1288 = n1287 ^ n1116 ;
  assign n1329 = n1328 ^ n1288 ;
  assign n1331 = n1010 & n1329 ;
  assign n1334 = n1331 ^ n1010 ;
  assign n1333 = n1009 & n1329 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1568 = n1567 ^ n1493 ;
  assign n1580 = n1579 ^ n1568 ;
  assign n1581 = n1580 ^ n1335 ;
  assign n1597 = n1596 ^ n1502 ;
  assign n1609 = n1608 ^ n1597 ;
  assign n1583 = n1041 & n1329 ;
  assign n1584 = n1583 ^ n1041 ;
  assign n1582 = n1040 & n1329 ;
  assign n1585 = n1584 ^ n1582 ;
  assign n1610 = n1609 ^ n1585 ;
  assign n1611 = n1581 & n1610 ;
  assign n1612 = n1611 ^ n1581 ;
  assign n1613 = n1612 ^ n1610 ;
  assign n1820 = n1335 & ~n1613 ;
  assign n1639 = n1049 & n1329 ;
  assign n1640 = n1639 ^ n1049 ;
  assign n1638 = n1077 & n1329 ;
  assign n1641 = n1640 ^ n1638 ;
  assign n1625 = n1624 ^ n1520 ;
  assign n1637 = n1636 ^ n1625 ;
  assign n1642 = n1641 ^ n1637 ;
  assign n1654 = n1653 ^ n1523 ;
  assign n1666 = n1665 ^ n1654 ;
  assign n1668 = n1080 & n1329 ;
  assign n1669 = n1668 ^ n1080 ;
  assign n1667 = n1108 & n1329 ;
  assign n1670 = n1669 ^ n1667 ;
  assign n1822 = n1666 & n1670 ;
  assign n1823 = n1822 ^ n1670 ;
  assign n1824 = n1642 & n1823 ;
  assign n1825 = n1824 ^ n1823 ;
  assign n1821 = ~n1637 & n1641 ;
  assign n1826 = n1825 ^ n1821 ;
  assign n1827 = n1820 & n1826 ;
  assign n1816 = n1585 & ~n1609 ;
  assign n1817 = ~n1581 & n1816 ;
  assign n1815 = n1335 & ~n1580 ;
  assign n1818 = n1817 ^ n1815 ;
  assign n1819 = n1335 & n1818 ;
  assign n1828 = n1827 ^ n1819 ;
  assign n2559 = n1828 ^ n1335 ;
  assign n1671 = n1670 ^ n1666 ;
  assign n1672 = n1642 & n1671 ;
  assign n1673 = n1672 ^ n1642 ;
  assign n1674 = n1673 ^ n1671 ;
  assign n1675 = n1613 & n1674 ;
  assign n1676 = n1675 ^ n1613 ;
  assign n1677 = n1676 ^ n1674 ;
  assign n1693 = n1692 ^ n1337 ;
  assign n1705 = n1704 ^ n1693 ;
  assign n1679 = n1124 & n1329 ;
  assign n1680 = n1679 ^ n1124 ;
  assign n1678 = n1152 & n1329 ;
  assign n1681 = n1680 ^ n1678 ;
  assign n1706 = n1705 ^ n1681 ;
  assign n1722 = n1721 ^ n1449 ;
  assign n1734 = n1733 ^ n1722 ;
  assign n1708 = n1155 & n1329 ;
  assign n1709 = n1708 ^ n1155 ;
  assign n1707 = n1183 & n1329 ;
  assign n1710 = n1709 ^ n1707 ;
  assign n1735 = n1734 ^ n1710 ;
  assign n1736 = n1706 & n1735 ;
  assign n1737 = n1736 ^ n1706 ;
  assign n1738 = n1737 ^ n1735 ;
  assign n1754 = n1753 ^ n1466 ;
  assign n1766 = n1765 ^ n1754 ;
  assign n1740 = n1200 & n1329 ;
  assign n1741 = n1740 ^ n1200 ;
  assign n1739 = n1289 & n1329 ;
  assign n1742 = n1741 ^ n1739 ;
  assign n1767 = n1766 ^ n1742 ;
  assign n1799 = n1205 & n1329 ;
  assign n1800 = n1799 ^ n1205 ;
  assign n1796 = n1318 & n1329 ;
  assign n1797 = n1796 ^ n1318 ;
  assign n1798 = n1797 ^ n1318 ;
  assign n1801 = n1800 ^ n1798 ;
  assign n1781 = n1780 ^ n1483 ;
  assign n1795 = n1794 ^ n1781 ;
  assign n1802 = n1801 ^ n1795 ;
  assign n1803 = n1767 & n1802 ;
  assign n1804 = n1803 ^ n1767 ;
  assign n1805 = n1804 ^ n1802 ;
  assign n1806 = n1738 & n1805 ;
  assign n1807 = n1806 ^ n1738 ;
  assign n1808 = n1807 ^ n1805 ;
  assign n1809 = n1677 & n1808 ;
  assign n1810 = n1809 ^ n1677 ;
  assign n1811 = n1810 ^ n1808 ;
  assign n1812 = n1335 & n1811 ;
  assign n1813 = n1812 ^ n1335 ;
  assign n1814 = n1813 ^ n1335 ;
  assign n2560 = n2559 ^ n1814 ;
  assign n1838 = n1795 & n1801 ;
  assign n1839 = n1838 ^ n1801 ;
  assign n1840 = n1767 & n1839 ;
  assign n1841 = n1840 ^ n1839 ;
  assign n1836 = n1742 & n1766 ;
  assign n1837 = n1836 ^ n1742 ;
  assign n1842 = n1841 ^ n1837 ;
  assign n1843 = n1738 & n1842 ;
  assign n1844 = n1843 ^ n1842 ;
  assign n1831 = n1710 & n1734 ;
  assign n1832 = n1831 ^ n1710 ;
  assign n1833 = n1706 & n1832 ;
  assign n1834 = n1833 ^ n1832 ;
  assign n1830 = n1681 & ~n1705 ;
  assign n1835 = n1834 ^ n1830 ;
  assign n1845 = n1844 ^ n1835 ;
  assign n1846 = n1335 & n1677 ;
  assign n1847 = n1846 ^ n1335 ;
  assign n1848 = n1845 & n1847 ;
  assign n2561 = n2560 ^ n1848 ;
  assign n1855 = n1580 & n1811 ;
  assign n1856 = n1855 ^ n1580 ;
  assign n1857 = n1856 ^ n1580 ;
  assign n1851 = n1580 & ~n1613 ;
  assign n1852 = n1826 & n1851 ;
  assign n1850 = n1580 & n1818 ;
  assign n1853 = n1852 ^ n1850 ;
  assign n2557 = n1857 ^ n1853 ;
  assign n1859 = n1580 & n1677 ;
  assign n1860 = n1859 ^ n1580 ;
  assign n1861 = n1845 & n1860 ;
  assign n2558 = n2557 ^ n1861 ;
  assign n2562 = n2561 ^ n2558 ;
  assign n2589 = n2588 ^ n2562 ;
  assign n2615 = n2367 & ~n2371 ;
  assign n2616 = n2422 & n2615 ;
  assign n2614 = n2367 & n2415 ;
  assign n2617 = n2616 ^ n2614 ;
  assign n2618 = n2617 ^ n2367 ;
  assign n2611 = n2367 & n2408 ;
  assign n2612 = n2611 ^ n2367 ;
  assign n2613 = n2612 ^ n2367 ;
  assign n2619 = n2618 ^ n2613 ;
  assign n2608 = n2367 & n2395 ;
  assign n2609 = n2608 ^ n2367 ;
  assign n2610 = n2350 & n2609 ;
  assign n2620 = n2619 ^ n2610 ;
  assign n2603 = n2361 & ~n2371 ;
  assign n2604 = n2422 & n2603 ;
  assign n2602 = n2361 & n2415 ;
  assign n2605 = n2604 ^ n2602 ;
  assign n2599 = n2361 & n2408 ;
  assign n2600 = n2599 ^ n2361 ;
  assign n2601 = n2600 ^ n2361 ;
  assign n2606 = n2605 ^ n2601 ;
  assign n2596 = n2361 & n2395 ;
  assign n2597 = n2596 ^ n2361 ;
  assign n2598 = n2350 & n2597 ;
  assign n2607 = n2606 ^ n2598 ;
  assign n2621 = n2620 ^ n2607 ;
  assign n1870 = n1585 & ~n1613 ;
  assign n1871 = n1826 & n1870 ;
  assign n1869 = n1585 & n1818 ;
  assign n1872 = n1871 ^ n1869 ;
  assign n2592 = n1872 ^ n1585 ;
  assign n1866 = n1585 & n1811 ;
  assign n1867 = n1866 ^ n1585 ;
  assign n1868 = n1867 ^ n1585 ;
  assign n2593 = n2592 ^ n1868 ;
  assign n1874 = n1585 & n1677 ;
  assign n1875 = n1874 ^ n1585 ;
  assign n1876 = n1845 & n1875 ;
  assign n2594 = n2593 ^ n1876 ;
  assign n1883 = n1609 & n1811 ;
  assign n1884 = n1883 ^ n1609 ;
  assign n1885 = n1884 ^ n1609 ;
  assign n1879 = n1609 & ~n1613 ;
  assign n1880 = n1826 & n1879 ;
  assign n1878 = n1609 & n1818 ;
  assign n1881 = n1880 ^ n1878 ;
  assign n2590 = n1885 ^ n1881 ;
  assign n1887 = n1609 & n1677 ;
  assign n1888 = n1887 ^ n1609 ;
  assign n1889 = n1845 & n1888 ;
  assign n2591 = n2590 ^ n1889 ;
  assign n2595 = n2594 ^ n2591 ;
  assign n2622 = n2621 ^ n2595 ;
  assign n2623 = n2589 & n2622 ;
  assign n2624 = n2623 ^ n2589 ;
  assign n2625 = n2624 ^ n2622 ;
  assign n2651 = ~n2371 & n2379 ;
  assign n2652 = n2422 & n2651 ;
  assign n2650 = n2379 & n2415 ;
  assign n2653 = n2652 ^ n2650 ;
  assign n2654 = n2653 ^ n2379 ;
  assign n2647 = n2379 & n2408 ;
  assign n2648 = n2647 ^ n2379 ;
  assign n2649 = n2648 ^ n2379 ;
  assign n2655 = n2654 ^ n2649 ;
  assign n2644 = n2379 & n2395 ;
  assign n2645 = n2644 ^ n2379 ;
  assign n2646 = n2350 & n2645 ;
  assign n2656 = n2655 ^ n2646 ;
  assign n2639 = ~n2371 & n2373 ;
  assign n2640 = n2422 & n2639 ;
  assign n2638 = n2373 & n2415 ;
  assign n2641 = n2640 ^ n2638 ;
  assign n2635 = n2373 & n2408 ;
  assign n2636 = n2635 ^ n2373 ;
  assign n2637 = n2636 ^ n2373 ;
  assign n2642 = n2641 ^ n2637 ;
  assign n2632 = n2373 & n2395 ;
  assign n2633 = n2632 ^ n2373 ;
  assign n2634 = n2350 & n2633 ;
  assign n2643 = n2642 ^ n2634 ;
  assign n2657 = n2656 ^ n2643 ;
  assign n1907 = ~n1613 & n1641 ;
  assign n1908 = n1826 & n1907 ;
  assign n1906 = n1641 & n1818 ;
  assign n1909 = n1908 ^ n1906 ;
  assign n2628 = n1909 ^ n1641 ;
  assign n1903 = n1641 & n1811 ;
  assign n1904 = n1903 ^ n1641 ;
  assign n1905 = n1904 ^ n1641 ;
  assign n2629 = n2628 ^ n1905 ;
  assign n1911 = n1641 & n1677 ;
  assign n1912 = n1911 ^ n1641 ;
  assign n1913 = n1845 & n1912 ;
  assign n2630 = n2629 ^ n1913 ;
  assign n1920 = n1637 & n1811 ;
  assign n1921 = n1920 ^ n1637 ;
  assign n1922 = n1921 ^ n1637 ;
  assign n1916 = ~n1613 & n1637 ;
  assign n1917 = n1826 & n1916 ;
  assign n1915 = n1637 & n1818 ;
  assign n1918 = n1917 ^ n1915 ;
  assign n2626 = n1922 ^ n1918 ;
  assign n1924 = n1637 & n1677 ;
  assign n1925 = n1924 ^ n1637 ;
  assign n1926 = n1845 & n1925 ;
  assign n2627 = n2626 ^ n1926 ;
  assign n2631 = n2630 ^ n2627 ;
  assign n2658 = n2657 ^ n2631 ;
  assign n1937 = ~n1613 & n1670 ;
  assign n1938 = n1826 & n1937 ;
  assign n1936 = n1670 & n1818 ;
  assign n1939 = n1938 ^ n1936 ;
  assign n2661 = n1939 ^ n1670 ;
  assign n1933 = n1670 & n1811 ;
  assign n1934 = n1933 ^ n1670 ;
  assign n1935 = n1934 ^ n1670 ;
  assign n2662 = n2661 ^ n1935 ;
  assign n1941 = n1670 & n1677 ;
  assign n1942 = n1941 ^ n1670 ;
  assign n1943 = n1845 & n1942 ;
  assign n2663 = n2662 ^ n1943 ;
  assign n1950 = n1666 & n1811 ;
  assign n1951 = n1950 ^ n1666 ;
  assign n1952 = n1951 ^ n1666 ;
  assign n1946 = ~n1613 & n1666 ;
  assign n1947 = n1826 & n1946 ;
  assign n1945 = n1666 & n1818 ;
  assign n1948 = n1947 ^ n1945 ;
  assign n2659 = n1952 ^ n1948 ;
  assign n1954 = n1666 & n1677 ;
  assign n1955 = n1954 ^ n1666 ;
  assign n1956 = n1845 & n1955 ;
  assign n2660 = n2659 ^ n1956 ;
  assign n2664 = n2663 ^ n2660 ;
  assign n2684 = ~n2371 & n2388 ;
  assign n2685 = n2422 & n2684 ;
  assign n2683 = n2388 & n2415 ;
  assign n2686 = n2685 ^ n2683 ;
  assign n2687 = n2686 ^ n2388 ;
  assign n2680 = n2388 & n2408 ;
  assign n2681 = n2680 ^ n2388 ;
  assign n2682 = n2681 ^ n2388 ;
  assign n2688 = n2687 ^ n2682 ;
  assign n2677 = n2388 & n2395 ;
  assign n2678 = n2677 ^ n2388 ;
  assign n2679 = n2350 & n2678 ;
  assign n2689 = n2688 ^ n2679 ;
  assign n2672 = ~n2371 & n2382 ;
  assign n2673 = n2422 & n2672 ;
  assign n2671 = n2382 & n2415 ;
  assign n2674 = n2673 ^ n2671 ;
  assign n2668 = n2382 & n2408 ;
  assign n2669 = n2668 ^ n2382 ;
  assign n2670 = n2669 ^ n2382 ;
  assign n2675 = n2674 ^ n2670 ;
  assign n2665 = n2382 & n2395 ;
  assign n2666 = n2665 ^ n2382 ;
  assign n2667 = n2350 & n2666 ;
  assign n2676 = n2675 ^ n2667 ;
  assign n2690 = n2689 ^ n2676 ;
  assign n2715 = n2664 & n2690 ;
  assign n2716 = n2715 ^ n2664 ;
  assign n2717 = n2658 & n2716 ;
  assign n2718 = n2717 ^ n2716 ;
  assign n2714 = n2631 & ~n2657 ;
  assign n2719 = n2718 ^ n2714 ;
  assign n2720 = n2625 & n2719 ;
  assign n2721 = n2720 ^ n2719 ;
  assign n2711 = n2595 & ~n2621 ;
  assign n2712 = ~n2589 & n2711 ;
  assign n2710 = n2562 & ~n2588 ;
  assign n2713 = n2712 ^ n2710 ;
  assign n2722 = n2721 ^ n2713 ;
  assign n2847 = n2588 & n2722 ;
  assign n2848 = n2847 ^ n2588 ;
  assign n2691 = n2690 ^ n2664 ;
  assign n2692 = n2658 & n2691 ;
  assign n2693 = n2692 ^ n2658 ;
  assign n2694 = n2693 ^ n2691 ;
  assign n2695 = n2625 & n2694 ;
  assign n2696 = n2695 ^ n2625 ;
  assign n2697 = n2696 ^ n2694 ;
  assign n2435 = n2304 & ~n2371 ;
  assign n2436 = n2422 & n2435 ;
  assign n2434 = n2304 & n2415 ;
  assign n2437 = n2436 ^ n2434 ;
  assign n2438 = n2437 ^ n2304 ;
  assign n2431 = n2304 & n2408 ;
  assign n2432 = n2431 ^ n2304 ;
  assign n2433 = n2432 ^ n2304 ;
  assign n2439 = n2438 ^ n2433 ;
  assign n2428 = n2304 & n2395 ;
  assign n2429 = n2428 ^ n2304 ;
  assign n2430 = n2350 & n2429 ;
  assign n2440 = n2439 ^ n2430 ;
  assign n2423 = n2195 & ~n2371 ;
  assign n2424 = n2422 & n2423 ;
  assign n2416 = n2195 & n2415 ;
  assign n2425 = n2424 ^ n2416 ;
  assign n2409 = n2195 & n2408 ;
  assign n2410 = n2409 ^ n2195 ;
  assign n2411 = n2410 ^ n2195 ;
  assign n2426 = n2425 ^ n2411 ;
  assign n2396 = n2195 & n2395 ;
  assign n2397 = n2396 ^ n2195 ;
  assign n2398 = n2350 & n2397 ;
  assign n2427 = n2426 ^ n2398 ;
  assign n2441 = n2440 ^ n2427 ;
  assign n1980 = ~n1613 & n1681 ;
  assign n1981 = n1826 & n1980 ;
  assign n1979 = n1681 & n1818 ;
  assign n1982 = n1981 ^ n1979 ;
  assign n2190 = n1982 ^ n1681 ;
  assign n1976 = n1681 & n1811 ;
  assign n1977 = n1976 ^ n1681 ;
  assign n1978 = n1977 ^ n1681 ;
  assign n2191 = n2190 ^ n1978 ;
  assign n1984 = n1677 & n1681 ;
  assign n1985 = n1984 ^ n1681 ;
  assign n1986 = n1845 & n1985 ;
  assign n2192 = n2191 ^ n1986 ;
  assign n1993 = n1705 & n1811 ;
  assign n1994 = n1993 ^ n1705 ;
  assign n1995 = n1994 ^ n1705 ;
  assign n1989 = ~n1613 & n1705 ;
  assign n1990 = n1826 & n1989 ;
  assign n1988 = n1705 & n1818 ;
  assign n1991 = n1990 ^ n1988 ;
  assign n2188 = n1995 ^ n1991 ;
  assign n1997 = n1677 & n1705 ;
  assign n1998 = n1997 ^ n1705 ;
  assign n1999 = n1845 & n1998 ;
  assign n2189 = n2188 ^ n1999 ;
  assign n2193 = n2192 ^ n2189 ;
  assign n2443 = n2441 ^ n2193 ;
  assign n2469 = n2314 & ~n2371 ;
  assign n2470 = n2422 & n2469 ;
  assign n2468 = n2314 & n2415 ;
  assign n2471 = n2470 ^ n2468 ;
  assign n2472 = n2471 ^ n2314 ;
  assign n2465 = n2314 & n2408 ;
  assign n2466 = n2465 ^ n2314 ;
  assign n2467 = n2466 ^ n2314 ;
  assign n2473 = n2472 ^ n2467 ;
  assign n2462 = n2314 & n2395 ;
  assign n2463 = n2462 ^ n2314 ;
  assign n2464 = n2350 & n2463 ;
  assign n2474 = n2473 ^ n2464 ;
  assign n2457 = n2308 & ~n2371 ;
  assign n2458 = n2422 & n2457 ;
  assign n2456 = n2308 & n2415 ;
  assign n2459 = n2458 ^ n2456 ;
  assign n2453 = n2308 & n2408 ;
  assign n2454 = n2453 ^ n2308 ;
  assign n2455 = n2454 ^ n2308 ;
  assign n2460 = n2459 ^ n2455 ;
  assign n2450 = n2308 & n2395 ;
  assign n2451 = n2450 ^ n2308 ;
  assign n2452 = n2350 & n2451 ;
  assign n2461 = n2460 ^ n2452 ;
  assign n2475 = n2474 ^ n2461 ;
  assign n2010 = ~n1613 & n1710 ;
  assign n2011 = n1826 & n2010 ;
  assign n2009 = n1710 & n1818 ;
  assign n2012 = n2011 ^ n2009 ;
  assign n2446 = n2012 ^ n1710 ;
  assign n2006 = n1710 & n1811 ;
  assign n2007 = n2006 ^ n1710 ;
  assign n2008 = n2007 ^ n1710 ;
  assign n2447 = n2446 ^ n2008 ;
  assign n2014 = n1677 & n1710 ;
  assign n2015 = n2014 ^ n1710 ;
  assign n2016 = n1845 & n2015 ;
  assign n2448 = n2447 ^ n2016 ;
  assign n2023 = n1734 & n1811 ;
  assign n2024 = n2023 ^ n1734 ;
  assign n2025 = n2024 ^ n1734 ;
  assign n2019 = ~n1613 & n1734 ;
  assign n2020 = n1826 & n2019 ;
  assign n2018 = n1734 & n1818 ;
  assign n2021 = n2020 ^ n2018 ;
  assign n2444 = n2025 ^ n2021 ;
  assign n2027 = n1677 & n1734 ;
  assign n2028 = n2027 ^ n1734 ;
  assign n2029 = n1845 & n2028 ;
  assign n2445 = n2444 ^ n2029 ;
  assign n2449 = n2448 ^ n2445 ;
  assign n2479 = n2475 ^ n2449 ;
  assign n2480 = n2443 & n2479 ;
  assign n2481 = n2480 ^ n2443 ;
  assign n2482 = n2481 ^ n2479 ;
  assign n2508 = n2331 & ~n2371 ;
  assign n2509 = n2422 & n2508 ;
  assign n2507 = n2331 & n2415 ;
  assign n2510 = n2509 ^ n2507 ;
  assign n2511 = n2510 ^ n2331 ;
  assign n2504 = n2331 & n2408 ;
  assign n2505 = n2504 ^ n2331 ;
  assign n2506 = n2505 ^ n2331 ;
  assign n2512 = n2511 ^ n2506 ;
  assign n2501 = n2331 & n2395 ;
  assign n2502 = n2501 ^ n2331 ;
  assign n2503 = n2350 & n2502 ;
  assign n2513 = n2512 ^ n2503 ;
  assign n2496 = n2325 & ~n2371 ;
  assign n2497 = n2422 & n2496 ;
  assign n2495 = n2325 & n2415 ;
  assign n2498 = n2497 ^ n2495 ;
  assign n2492 = n2325 & n2408 ;
  assign n2493 = n2492 ^ n2325 ;
  assign n2494 = n2493 ^ n2325 ;
  assign n2499 = n2498 ^ n2494 ;
  assign n2489 = n2325 & n2395 ;
  assign n2490 = n2489 ^ n2325 ;
  assign n2491 = n2350 & n2490 ;
  assign n2500 = n2499 ^ n2491 ;
  assign n2514 = n2513 ^ n2500 ;
  assign n2094 = ~n1613 & n1742 ;
  assign n2095 = n1826 & n2094 ;
  assign n2093 = n1742 & n1818 ;
  assign n2096 = n2095 ^ n2093 ;
  assign n2485 = n2096 ^ n1742 ;
  assign n2089 = n1742 & n1811 ;
  assign n2090 = n2089 ^ n1742 ;
  assign n2091 = n2090 ^ n1742 ;
  assign n2486 = n2485 ^ n2091 ;
  assign n2084 = n1677 & n1742 ;
  assign n2137 = n2084 ^ n1742 ;
  assign n2138 = n1845 & n2137 ;
  assign n2487 = n2486 ^ n2138 ;
  assign n2111 = ~n1613 & n1766 ;
  assign n2112 = n1826 & n2111 ;
  assign n2110 = n1766 & n1818 ;
  assign n2113 = n2112 ^ n2110 ;
  assign n2106 = n1766 & n1811 ;
  assign n2107 = n2106 ^ n1766 ;
  assign n2108 = n2107 ^ n1766 ;
  assign n2483 = n2113 ^ n2108 ;
  assign n2101 = n1677 & n1766 ;
  assign n2142 = n2101 ^ n1766 ;
  assign n2143 = n1845 & n2142 ;
  assign n2484 = n2483 ^ n2143 ;
  assign n2488 = n2487 ^ n2484 ;
  assign n2516 = n2514 ^ n2488 ;
  assign n2543 = n2342 & ~n2371 ;
  assign n2544 = n2422 & n2543 ;
  assign n2542 = n2342 & ~n2415 ;
  assign n2545 = n2544 ^ n2542 ;
  assign n2539 = n2342 & n2408 ;
  assign n2540 = n2539 ^ n2342 ;
  assign n2541 = n2540 ^ n2342 ;
  assign n2546 = n2545 ^ n2541 ;
  assign n2536 = n2342 & n2395 ;
  assign n2537 = n2536 ^ n2342 ;
  assign n2538 = n2350 & n2537 ;
  assign n2547 = n2546 ^ n2538 ;
  assign n2530 = n2336 & ~n2371 ;
  assign n2531 = n2422 & n2530 ;
  assign n2529 = n2336 & ~n2415 ;
  assign n2532 = n2531 ^ n2529 ;
  assign n2526 = n2336 & n2408 ;
  assign n2527 = n2526 ^ n2336 ;
  assign n2528 = n2527 ^ n2336 ;
  assign n2533 = n2532 ^ n2528 ;
  assign n2523 = n2336 & n2395 ;
  assign n2524 = n2523 ^ n2336 ;
  assign n2525 = n2350 & n2524 ;
  assign n2534 = n2533 ^ n2525 ;
  assign n2535 = n2534 ^ n2336 ;
  assign n2548 = n2547 ^ n2535 ;
  assign n2518 = n1801 & ~n1818 ;
  assign n2148 = ~n1613 & n1801 ;
  assign n2149 = n1826 & n2148 ;
  assign n2519 = n2518 ^ n2149 ;
  assign n2151 = n1801 & n1811 ;
  assign n2152 = n2151 ^ n1801 ;
  assign n2153 = n2152 ^ n1801 ;
  assign n2520 = n2519 ^ n2153 ;
  assign n2155 = n1677 & n1801 ;
  assign n2156 = n2155 ^ n1801 ;
  assign n2157 = n1845 & n2156 ;
  assign n2521 = n2520 ^ n2157 ;
  assign n2166 = ~n1613 & n1795 ;
  assign n2167 = n1826 & n2166 ;
  assign n2165 = n1795 & ~n1818 ;
  assign n2168 = n2167 ^ n2165 ;
  assign n2162 = n1795 & n1811 ;
  assign n2163 = n2162 ^ n1795 ;
  assign n2164 = n2163 ^ n1795 ;
  assign n2169 = n2168 ^ n2164 ;
  assign n2159 = n1677 & n1795 ;
  assign n2160 = n2159 ^ n1795 ;
  assign n2161 = n1845 & n2160 ;
  assign n2170 = n2169 ^ n2161 ;
  assign n2517 = n2170 ^ n1795 ;
  assign n2522 = n2521 ^ n2517 ;
  assign n2700 = n2548 ^ n2522 ;
  assign n2701 = n2516 & n2700 ;
  assign n2702 = n2701 ^ n2516 ;
  assign n2703 = n2702 ^ n2700 ;
  assign n2704 = n2482 & n2703 ;
  assign n2705 = n2704 ^ n2482 ;
  assign n2706 = n2705 ^ n2703 ;
  assign n2707 = ~n2697 & ~n2706 ;
  assign n2845 = n2588 & n2707 ;
  assign n2846 = n2845 ^ n2588 ;
  assign n2849 = n2848 ^ n2846 ;
  assign n2549 = n2522 & n2548 ;
  assign n2550 = n2549 ^ n2522 ;
  assign n2551 = n2516 & n2550 ;
  assign n2552 = n2551 ^ n2550 ;
  assign n2515 = n2488 & ~n2514 ;
  assign n2553 = n2552 ^ n2515 ;
  assign n2554 = n2482 & n2553 ;
  assign n2555 = n2554 ^ n2553 ;
  assign n2476 = n2449 & ~n2475 ;
  assign n2477 = ~n2443 & n2476 ;
  assign n2442 = n2193 & ~n2441 ;
  assign n2478 = n2477 ^ n2442 ;
  assign n2556 = n2555 ^ n2478 ;
  assign n2843 = n2588 & ~n2697 ;
  assign n2844 = n2556 & n2843 ;
  assign n2850 = n2849 ^ n2844 ;
  assign n2838 = n2562 & n2722 ;
  assign n2839 = n2838 ^ n2562 ;
  assign n2836 = n2562 & n2707 ;
  assign n2837 = n2836 ^ n2562 ;
  assign n2840 = n2839 ^ n2837 ;
  assign n2834 = n2562 & ~n2697 ;
  assign n2835 = n2556 & n2834 ;
  assign n2841 = n2840 ^ n2835 ;
  assign n2842 = n2841 ^ n2562 ;
  assign n2851 = n2850 ^ n2842 ;
  assign n1330 = n1009 & ~n1329 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1854 = n1853 ^ n1580 ;
  assign n1858 = n1857 ^ n1854 ;
  assign n1862 = n1861 ^ n1858 ;
  assign n1829 = n1828 ^ n1814 ;
  assign n1849 = n1848 ^ n1829 ;
  assign n1863 = n1862 ^ n1849 ;
  assign n1865 = n1863 ^ n1332 ;
  assign n1892 = n1040 & ~n1329 ;
  assign n1893 = n1892 ^ n1583 ;
  assign n1882 = n1881 ^ n1609 ;
  assign n1886 = n1885 ^ n1882 ;
  assign n1890 = n1889 ^ n1886 ;
  assign n1873 = n1872 ^ n1868 ;
  assign n1877 = n1876 ^ n1873 ;
  assign n1891 = n1890 ^ n1877 ;
  assign n1897 = n1893 ^ n1891 ;
  assign n1898 = n1865 & n1897 ;
  assign n1899 = n1898 ^ n1865 ;
  assign n1900 = n1899 ^ n1897 ;
  assign n1919 = n1918 ^ n1637 ;
  assign n1923 = n1922 ^ n1919 ;
  assign n1927 = n1926 ^ n1923 ;
  assign n1910 = n1909 ^ n1905 ;
  assign n1914 = n1913 ^ n1910 ;
  assign n1928 = n1927 ^ n1914 ;
  assign n1901 = n1077 & ~n1329 ;
  assign n1902 = n1901 ^ n1639 ;
  assign n1930 = n1928 ^ n1902 ;
  assign n1949 = n1948 ^ n1666 ;
  assign n1953 = n1952 ^ n1949 ;
  assign n1957 = n1956 ^ n1953 ;
  assign n1940 = n1939 ^ n1935 ;
  assign n1944 = n1943 ^ n1940 ;
  assign n1958 = n1957 ^ n1944 ;
  assign n1931 = n1108 & ~n1329 ;
  assign n1932 = n1931 ^ n1668 ;
  assign n1967 = n1958 ^ n1932 ;
  assign n1968 = n1930 & n1967 ;
  assign n1969 = n1968 ^ n1930 ;
  assign n1970 = n1969 ^ n1967 ;
  assign n1971 = n1900 & n1970 ;
  assign n1972 = n1971 ^ n1900 ;
  assign n1973 = n1972 ^ n1970 ;
  assign n1992 = n1991 ^ n1705 ;
  assign n1996 = n1995 ^ n1992 ;
  assign n2000 = n1999 ^ n1996 ;
  assign n1983 = n1982 ^ n1978 ;
  assign n1987 = n1986 ^ n1983 ;
  assign n2001 = n2000 ^ n1987 ;
  assign n1974 = n1152 & ~n1329 ;
  assign n1975 = n1974 ^ n1679 ;
  assign n2003 = n2001 ^ n1975 ;
  assign n2022 = n2021 ^ n1734 ;
  assign n2026 = n2025 ^ n2022 ;
  assign n2030 = n2029 ^ n2026 ;
  assign n2013 = n2012 ^ n2008 ;
  assign n2017 = n2016 ^ n2013 ;
  assign n2031 = n2030 ^ n2017 ;
  assign n2004 = n1183 & ~n1329 ;
  assign n2005 = n2004 ^ n1708 ;
  assign n2037 = n2031 ^ n2005 ;
  assign n2038 = n2003 & n2037 ;
  assign n2039 = n2038 ^ n2003 ;
  assign n2040 = n2039 ^ n2037 ;
  assign n2140 = n2113 ^ n1766 ;
  assign n2141 = n2140 ^ n2108 ;
  assign n2144 = n2143 ^ n2141 ;
  assign n2136 = n2096 ^ n2091 ;
  assign n2139 = n2138 ^ n2136 ;
  assign n2145 = n2144 ^ n2139 ;
  assign n2048 = n1289 & ~n1329 ;
  assign n2049 = n2048 ^ n1740 ;
  assign n2146 = n2145 ^ n2049 ;
  assign n2147 = n1801 & n1818 ;
  assign n2150 = n2149 ^ n2147 ;
  assign n2154 = n2153 ^ n2150 ;
  assign n2158 = n2157 ^ n2154 ;
  assign n2171 = n2170 ^ n2158 ;
  assign n2054 = n1799 ^ n1797 ;
  assign n2172 = n2171 ^ n2054 ;
  assign n2173 = n2146 & n2172 ;
  assign n2174 = n2173 ^ n2146 ;
  assign n2175 = n2174 ^ n2172 ;
  assign n2176 = n2040 & n2175 ;
  assign n2177 = n2176 ^ n2040 ;
  assign n2178 = n2177 ^ n2175 ;
  assign n2179 = ~n1973 & ~n2178 ;
  assign n2122 = ~n1766 & n2049 ;
  assign n2126 = n1811 & n2122 ;
  assign n2043 = n1613 & n1826 ;
  assign n2044 = n2043 ^ n1826 ;
  assign n2045 = n2044 ^ n1818 ;
  assign n2125 = ~n2045 & n2122 ;
  assign n2127 = n2126 ^ n2125 ;
  assign n2123 = ~n1677 & n2122 ;
  assign n2124 = n1845 & n2123 ;
  assign n2128 = n2127 ^ n2124 ;
  assign n2069 = ~n1801 & n2054 ;
  assign n2077 = ~n1613 & n2069 ;
  assign n2078 = n1826 & n2077 ;
  assign n2076 = n1818 & n2069 ;
  assign n2079 = n2078 ^ n2076 ;
  assign n2073 = n1811 & n2069 ;
  assign n2074 = n2073 ^ n2069 ;
  assign n2075 = n2074 ^ n2069 ;
  assign n2080 = n2079 ^ n2075 ;
  assign n2070 = n1677 & n2069 ;
  assign n2071 = n2070 ^ n2069 ;
  assign n2072 = n1845 & n2071 ;
  assign n2081 = n2080 ^ n2072 ;
  assign n2055 = ~n1795 & n2054 ;
  assign n2063 = ~n1613 & n2055 ;
  assign n2064 = n1826 & n2063 ;
  assign n2062 = n1818 & n2055 ;
  assign n2065 = n2064 ^ n2062 ;
  assign n2066 = n2065 ^ n2055 ;
  assign n2059 = n1811 & n2055 ;
  assign n2060 = n2059 ^ n2055 ;
  assign n2061 = n2060 ^ n2055 ;
  assign n2067 = n2066 ^ n2061 ;
  assign n2056 = n1677 & n2055 ;
  assign n2057 = n2056 ^ n2055 ;
  assign n2058 = n1845 & n2057 ;
  assign n2068 = n2067 ^ n2058 ;
  assign n2082 = n2081 ^ n2068 ;
  assign n2114 = n2113 ^ n2045 ;
  assign n2115 = n2114 ^ n1766 ;
  assign n2109 = n2108 ^ n1811 ;
  assign n2116 = n2115 ^ n2109 ;
  assign n2102 = n2101 ^ n1677 ;
  assign n2103 = n2102 ^ n1766 ;
  assign n2104 = n1845 & n2103 ;
  assign n2105 = n2104 ^ n1845 ;
  assign n2117 = n2116 ^ n2105 ;
  assign n2118 = n2082 & n2117 ;
  assign n2119 = n2118 ^ n2082 ;
  assign n2097 = n2096 ^ n2045 ;
  assign n2092 = n2091 ^ n1811 ;
  assign n2098 = n2097 ^ n2092 ;
  assign n2085 = n2084 ^ n1677 ;
  assign n2086 = n2085 ^ n1742 ;
  assign n2087 = n1845 & n2086 ;
  assign n2088 = n2087 ^ n1845 ;
  assign n2099 = n2098 ^ n2088 ;
  assign n2100 = n2082 & n2099 ;
  assign n2120 = n2119 ^ n2100 ;
  assign n2083 = n2049 & n2082 ;
  assign n2121 = n2120 ^ n2083 ;
  assign n2129 = n2128 ^ n2121 ;
  assign n2041 = n1677 & n1845 ;
  assign n2042 = n2041 ^ n1845 ;
  assign n2046 = n2045 ^ n2042 ;
  assign n2047 = n2046 ^ n1811 ;
  assign n2050 = ~n1742 & n2049 ;
  assign n2051 = n2047 & n2050 ;
  assign n2052 = n2051 ^ n2050 ;
  assign n2053 = n2052 ^ n2050 ;
  assign n2130 = n2129 ^ n2053 ;
  assign n2131 = n2040 & n2130 ;
  assign n2132 = n2131 ^ n2130 ;
  assign n2032 = n2005 & n2031 ;
  assign n2033 = n2032 ^ n2005 ;
  assign n2034 = n2003 & n2033 ;
  assign n2035 = n2034 ^ n2033 ;
  assign n2002 = n1975 & ~n2001 ;
  assign n2036 = n2035 ^ n2002 ;
  assign n2133 = n2132 ^ n2036 ;
  assign n2134 = ~n1973 & n2133 ;
  assign n1959 = n1932 & n1958 ;
  assign n1960 = n1959 ^ n1932 ;
  assign n1961 = n1930 & n1960 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1929 = n1902 & ~n1928 ;
  assign n1963 = n1962 ^ n1929 ;
  assign n1964 = n1900 & n1963 ;
  assign n1965 = n1964 ^ n1963 ;
  assign n1894 = ~n1891 & n1893 ;
  assign n1895 = ~n1865 & n1894 ;
  assign n1864 = n1332 & ~n1863 ;
  assign n1896 = n1895 ^ n1864 ;
  assign n1966 = n1965 ^ n1896 ;
  assign n2135 = n2134 ^ n1966 ;
  assign n2180 = n2179 ^ n2135 ;
  assign n2832 = n1332 & n2180 ;
  assign n2182 = n1863 & n2180 ;
  assign n2831 = n2182 ^ n1863 ;
  assign n2833 = n2832 ^ n2831 ;
  assign n2852 = n2851 ^ n2833 ;
  assign n2870 = n2621 & n2722 ;
  assign n2871 = n2870 ^ n2621 ;
  assign n2868 = n2621 & n2707 ;
  assign n2869 = n2868 ^ n2621 ;
  assign n2872 = n2871 ^ n2869 ;
  assign n2866 = n2621 & ~n2697 ;
  assign n2867 = n2556 & n2866 ;
  assign n2873 = n2872 ^ n2867 ;
  assign n2861 = n2595 & n2722 ;
  assign n2862 = n2861 ^ n2595 ;
  assign n2859 = n2595 & n2707 ;
  assign n2860 = n2859 ^ n2595 ;
  assign n2863 = n2862 ^ n2860 ;
  assign n2857 = n2595 & ~n2697 ;
  assign n2858 = n2556 & n2857 ;
  assign n2864 = n2863 ^ n2858 ;
  assign n2865 = n2864 ^ n2595 ;
  assign n2874 = n2873 ^ n2865 ;
  assign n2855 = n1893 & n2180 ;
  assign n2853 = n1891 & n2180 ;
  assign n2854 = n2853 ^ n1891 ;
  assign n2856 = n2855 ^ n2854 ;
  assign n2875 = n2874 ^ n2856 ;
  assign n2876 = n2852 & n2875 ;
  assign n2877 = n2876 ^ n2852 ;
  assign n2878 = n2877 ^ n2875 ;
  assign n2896 = n2657 & n2722 ;
  assign n2897 = n2896 ^ n2657 ;
  assign n2894 = n2657 & n2707 ;
  assign n2895 = n2894 ^ n2657 ;
  assign n2898 = n2897 ^ n2895 ;
  assign n2892 = n2657 & ~n2697 ;
  assign n2893 = n2556 & n2892 ;
  assign n2899 = n2898 ^ n2893 ;
  assign n2887 = n2631 & n2722 ;
  assign n2888 = n2887 ^ n2631 ;
  assign n2885 = n2631 & n2707 ;
  assign n2886 = n2885 ^ n2631 ;
  assign n2889 = n2888 ^ n2886 ;
  assign n2883 = n2631 & ~n2697 ;
  assign n2884 = n2556 & n2883 ;
  assign n2890 = n2889 ^ n2884 ;
  assign n2891 = n2890 ^ n2631 ;
  assign n2900 = n2899 ^ n2891 ;
  assign n2881 = n1902 & n2180 ;
  assign n2879 = n1928 & n2180 ;
  assign n2880 = n2879 ^ n1928 ;
  assign n2882 = n2881 ^ n2880 ;
  assign n2901 = n2900 ^ n2882 ;
  assign n2904 = n1932 & n2180 ;
  assign n2902 = n1958 & n2180 ;
  assign n2903 = n2902 ^ n1958 ;
  assign n2905 = n2904 ^ n2903 ;
  assign n2919 = n2690 & n2722 ;
  assign n2920 = n2919 ^ n2690 ;
  assign n2917 = n2690 & n2707 ;
  assign n2918 = n2917 ^ n2690 ;
  assign n2921 = n2920 ^ n2918 ;
  assign n2915 = n2690 & ~n2697 ;
  assign n2916 = n2556 & n2915 ;
  assign n2922 = n2921 ^ n2916 ;
  assign n2910 = n2664 & n2722 ;
  assign n2911 = n2910 ^ n2664 ;
  assign n2908 = n2664 & n2707 ;
  assign n2909 = n2908 ^ n2664 ;
  assign n2912 = n2911 ^ n2909 ;
  assign n2906 = n2664 & ~n2697 ;
  assign n2907 = n2556 & n2906 ;
  assign n2913 = n2912 ^ n2907 ;
  assign n2914 = n2913 ^ n2664 ;
  assign n2923 = n2922 ^ n2914 ;
  assign n2948 = n2905 & n2923 ;
  assign n2949 = n2948 ^ n2905 ;
  assign n2950 = n2901 & n2949 ;
  assign n2951 = n2950 ^ n2949 ;
  assign n2947 = n2882 & ~n2900 ;
  assign n2952 = n2951 ^ n2947 ;
  assign n2953 = n2878 & n2952 ;
  assign n2954 = n2953 ^ n2952 ;
  assign n2944 = n2856 & ~n2874 ;
  assign n2945 = ~n2852 & n2944 ;
  assign n2943 = n2833 & ~n2851 ;
  assign n2946 = n2945 ^ n2943 ;
  assign n2955 = n2954 ^ n2946 ;
  assign n2965 = n2851 & n2955 ;
  assign n2966 = n2965 ^ n2851 ;
  assign n2924 = n2923 ^ n2905 ;
  assign n2925 = n2901 & n2924 ;
  assign n2926 = n2925 ^ n2901 ;
  assign n2927 = n2926 ^ n2924 ;
  assign n2928 = n2878 & n2927 ;
  assign n2929 = n2928 ^ n2878 ;
  assign n2930 = n2929 ^ n2927 ;
  assign n2732 = n2441 & n2722 ;
  assign n2733 = n2732 ^ n2441 ;
  assign n2730 = n2441 & n2707 ;
  assign n2731 = n2730 ^ n2441 ;
  assign n2734 = n2733 ^ n2731 ;
  assign n2728 = n2441 & ~n2697 ;
  assign n2729 = n2556 & n2728 ;
  assign n2735 = n2734 ^ n2729 ;
  assign n2723 = n2193 & n2722 ;
  assign n2724 = n2723 ^ n2193 ;
  assign n2708 = n2193 & n2707 ;
  assign n2709 = n2708 ^ n2193 ;
  assign n2725 = n2724 ^ n2709 ;
  assign n2698 = n2193 & ~n2697 ;
  assign n2699 = n2556 & n2698 ;
  assign n2726 = n2725 ^ n2699 ;
  assign n2727 = n2726 ^ n2193 ;
  assign n2736 = n2735 ^ n2727 ;
  assign n2186 = n1975 & n2180 ;
  assign n2184 = n2001 & n2180 ;
  assign n2185 = n2184 ^ n2001 ;
  assign n2187 = n2186 ^ n2185 ;
  assign n2738 = n2736 ^ n2187 ;
  assign n2756 = n2475 & n2722 ;
  assign n2757 = n2756 ^ n2475 ;
  assign n2754 = n2475 & n2707 ;
  assign n2755 = n2754 ^ n2475 ;
  assign n2758 = n2757 ^ n2755 ;
  assign n2752 = n2475 & ~n2697 ;
  assign n2753 = n2556 & n2752 ;
  assign n2759 = n2758 ^ n2753 ;
  assign n2747 = n2449 & n2722 ;
  assign n2748 = n2747 ^ n2449 ;
  assign n2745 = n2449 & n2707 ;
  assign n2746 = n2745 ^ n2449 ;
  assign n2749 = n2748 ^ n2746 ;
  assign n2743 = n2449 & ~n2697 ;
  assign n2744 = n2556 & n2743 ;
  assign n2750 = n2749 ^ n2744 ;
  assign n2751 = n2750 ^ n2449 ;
  assign n2760 = n2759 ^ n2751 ;
  assign n2741 = n2005 & n2180 ;
  assign n2739 = n2031 & n2180 ;
  assign n2740 = n2739 ^ n2031 ;
  assign n2742 = n2741 ^ n2740 ;
  assign n2766 = n2760 ^ n2742 ;
  assign n2767 = n2738 & n2766 ;
  assign n2768 = n2767 ^ n2738 ;
  assign n2769 = n2768 ^ n2766 ;
  assign n2787 = n2514 & n2722 ;
  assign n2788 = n2787 ^ n2514 ;
  assign n2785 = n2514 & n2707 ;
  assign n2786 = n2785 ^ n2514 ;
  assign n2789 = n2788 ^ n2786 ;
  assign n2783 = n2514 & ~n2697 ;
  assign n2784 = n2556 & n2783 ;
  assign n2790 = n2789 ^ n2784 ;
  assign n2778 = n2488 & n2722 ;
  assign n2779 = n2778 ^ n2488 ;
  assign n2776 = n2488 & n2707 ;
  assign n2777 = n2776 ^ n2488 ;
  assign n2780 = n2779 ^ n2777 ;
  assign n2774 = n2488 & ~n2697 ;
  assign n2775 = n2556 & n2774 ;
  assign n2781 = n2780 ^ n2775 ;
  assign n2782 = n2781 ^ n2488 ;
  assign n2791 = n2790 ^ n2782 ;
  assign n2772 = n2049 & n2180 ;
  assign n2770 = n2145 & n2180 ;
  assign n2771 = n2770 ^ n2145 ;
  assign n2773 = n2772 ^ n2771 ;
  assign n2794 = n2791 ^ n2773 ;
  assign n2816 = n2548 & ~n2625 ;
  assign n2817 = n2719 & n2816 ;
  assign n2815 = n2548 & n2713 ;
  assign n2818 = n2817 ^ n2815 ;
  assign n2819 = n2818 ^ n2548 ;
  assign n2813 = n2548 & n2707 ;
  assign n2814 = n2813 ^ n2548 ;
  assign n2820 = n2819 ^ n2814 ;
  assign n2811 = n2548 & ~n2697 ;
  assign n2812 = n2556 & n2811 ;
  assign n2821 = n2820 ^ n2812 ;
  assign n2804 = n2522 & ~n2625 ;
  assign n2805 = n2719 & n2804 ;
  assign n2803 = n2522 & n2713 ;
  assign n2806 = n2805 ^ n2803 ;
  assign n2807 = n2806 ^ n2522 ;
  assign n2801 = n2522 & n2707 ;
  assign n2802 = n2801 ^ n2522 ;
  assign n2808 = n2807 ^ n2802 ;
  assign n2799 = n2522 & ~n2697 ;
  assign n2800 = n2556 & n2799 ;
  assign n2809 = n2808 ^ n2800 ;
  assign n2810 = n2809 ^ n2522 ;
  assign n2822 = n2821 ^ n2810 ;
  assign n2797 = n2054 & n2180 ;
  assign n2795 = n2171 & n2180 ;
  assign n2796 = n2795 ^ n2171 ;
  assign n2798 = n2797 ^ n2796 ;
  assign n2933 = n2822 ^ n2798 ;
  assign n2934 = n2794 & n2933 ;
  assign n2935 = n2934 ^ n2794 ;
  assign n2936 = n2935 ^ n2933 ;
  assign n2937 = n2769 & n2936 ;
  assign n2938 = n2937 ^ n2769 ;
  assign n2939 = n2938 ^ n2936 ;
  assign n2940 = ~n2930 & ~n2939 ;
  assign n2963 = n2851 & n2940 ;
  assign n2964 = n2963 ^ n2851 ;
  assign n2967 = n2966 ^ n2964 ;
  assign n2823 = n2798 & n2822 ;
  assign n2824 = n2823 ^ n2798 ;
  assign n2825 = n2794 & n2824 ;
  assign n2826 = n2825 ^ n2824 ;
  assign n2792 = n2773 & n2791 ;
  assign n2793 = n2792 ^ n2773 ;
  assign n2827 = n2826 ^ n2793 ;
  assign n2828 = n2769 & n2827 ;
  assign n2829 = n2828 ^ n2827 ;
  assign n2761 = n2742 & n2760 ;
  assign n2762 = n2761 ^ n2742 ;
  assign n2763 = n2738 & n2762 ;
  assign n2764 = n2763 ^ n2762 ;
  assign n2737 = n2187 & ~n2736 ;
  assign n2765 = n2764 ^ n2737 ;
  assign n2830 = n2829 ^ n2765 ;
  assign n2961 = n2851 & ~n2930 ;
  assign n2962 = n2830 & n2961 ;
  assign n2968 = n2967 ^ n2962 ;
  assign n2956 = n2833 & n2955 ;
  assign n2957 = n2956 ^ n2833 ;
  assign n2941 = n2833 & n2940 ;
  assign n2942 = n2941 ^ n2833 ;
  assign n2958 = n2957 ^ n2942 ;
  assign n2931 = n2833 & ~n2930 ;
  assign n2932 = n2830 & n2931 ;
  assign n2959 = n2958 ^ n2932 ;
  assign n2960 = n2959 ^ n2833 ;
  assign n2969 = n2968 ^ n2960 ;
  assign n2181 = n1332 & ~n2180 ;
  assign n2183 = n2182 ^ n2181 ;
  assign n2994 = n2969 ^ n2183 ;
  assign n2989 = n1893 & ~n2180 ;
  assign n2990 = n2989 ^ n2853 ;
  assign n2984 = n2874 & n2955 ;
  assign n2985 = n2984 ^ n2874 ;
  assign n2982 = n2874 & n2940 ;
  assign n2983 = n2982 ^ n2874 ;
  assign n2986 = n2985 ^ n2983 ;
  assign n2980 = n2874 & ~n2930 ;
  assign n2981 = n2830 & n2980 ;
  assign n2987 = n2986 ^ n2981 ;
  assign n2975 = n2856 & n2955 ;
  assign n2976 = n2975 ^ n2856 ;
  assign n2973 = n2856 & n2940 ;
  assign n2974 = n2973 ^ n2856 ;
  assign n2977 = n2976 ^ n2974 ;
  assign n2971 = n2856 & ~n2930 ;
  assign n2972 = n2830 & n2971 ;
  assign n2978 = n2977 ^ n2972 ;
  assign n2979 = n2978 ^ n2856 ;
  assign n2988 = n2987 ^ n2979 ;
  assign n2995 = n2990 ^ n2988 ;
  assign n2996 = n2994 & n2995 ;
  assign n2997 = n2996 ^ n2994 ;
  assign n2998 = n2997 ^ n2995 ;
  assign n3014 = n2900 & n2955 ;
  assign n3015 = n3014 ^ n2900 ;
  assign n3012 = n2900 & n2940 ;
  assign n3013 = n3012 ^ n2900 ;
  assign n3016 = n3015 ^ n3013 ;
  assign n3010 = n2900 & ~n2930 ;
  assign n3011 = n2830 & n3010 ;
  assign n3017 = n3016 ^ n3011 ;
  assign n3005 = n2882 & n2955 ;
  assign n3006 = n3005 ^ n2882 ;
  assign n3003 = n2882 & n2940 ;
  assign n3004 = n3003 ^ n2882 ;
  assign n3007 = n3006 ^ n3004 ;
  assign n3001 = n2882 & ~n2930 ;
  assign n3002 = n2830 & n3001 ;
  assign n3008 = n3007 ^ n3002 ;
  assign n3009 = n3008 ^ n2882 ;
  assign n3018 = n3017 ^ n3009 ;
  assign n2999 = n1902 & ~n2180 ;
  assign n3000 = n2999 ^ n2879 ;
  assign n3020 = n3018 ^ n3000 ;
  assign n3055 = n2923 & n2955 ;
  assign n3056 = n3055 ^ n2923 ;
  assign n3053 = n2923 & n2940 ;
  assign n3054 = n3053 ^ n2923 ;
  assign n3057 = n3056 ^ n3054 ;
  assign n3051 = n2923 & ~n2930 ;
  assign n3052 = n2830 & n3051 ;
  assign n3058 = n3057 ^ n3052 ;
  assign n3046 = n2905 & n2955 ;
  assign n3047 = n3046 ^ n2905 ;
  assign n3044 = n2905 & n2940 ;
  assign n3045 = n3044 ^ n2905 ;
  assign n3048 = n3047 ^ n3045 ;
  assign n3042 = n2905 & ~n2930 ;
  assign n3043 = n2830 & n3042 ;
  assign n3049 = n3048 ^ n3043 ;
  assign n3050 = n3049 ^ n2905 ;
  assign n3059 = n3058 ^ n3050 ;
  assign n3024 = n1932 & ~n2180 ;
  assign n3025 = n3024 ^ n2902 ;
  assign n3060 = n3059 ^ n3025 ;
  assign n3061 = n3020 & n3060 ;
  assign n3062 = n3061 ^ n3020 ;
  assign n3063 = n3062 ^ n3060 ;
  assign n3064 = n2998 & n3063 ;
  assign n3065 = n3064 ^ n2998 ;
  assign n3066 = n3065 ^ n3063 ;
  assign n3082 = n2736 & n2955 ;
  assign n3083 = n3082 ^ n2736 ;
  assign n3080 = n2736 & n2940 ;
  assign n3081 = n3080 ^ n2736 ;
  assign n3084 = n3083 ^ n3081 ;
  assign n3078 = n2736 & ~n2930 ;
  assign n3079 = n2830 & n3078 ;
  assign n3085 = n3084 ^ n3079 ;
  assign n3073 = n2187 & n2955 ;
  assign n3074 = n3073 ^ n2187 ;
  assign n3071 = n2187 & n2940 ;
  assign n3072 = n3071 ^ n2187 ;
  assign n3075 = n3074 ^ n3072 ;
  assign n3069 = n2187 & ~n2930 ;
  assign n3070 = n2830 & n3069 ;
  assign n3076 = n3075 ^ n3070 ;
  assign n3077 = n3076 ^ n2187 ;
  assign n3086 = n3085 ^ n3077 ;
  assign n3067 = n1975 & ~n2180 ;
  assign n3068 = n3067 ^ n2184 ;
  assign n3088 = n3086 ^ n3068 ;
  assign n3114 = n2760 & n2955 ;
  assign n3115 = n3114 ^ n2760 ;
  assign n3112 = n2760 & n2940 ;
  assign n3113 = n3112 ^ n2760 ;
  assign n3116 = n3115 ^ n3113 ;
  assign n3110 = n2760 & ~n2930 ;
  assign n3111 = n2830 & n3110 ;
  assign n3117 = n3116 ^ n3111 ;
  assign n3105 = n2742 & n2955 ;
  assign n3106 = n3105 ^ n2742 ;
  assign n3103 = n2742 & n2940 ;
  assign n3104 = n3103 ^ n2742 ;
  assign n3107 = n3106 ^ n3104 ;
  assign n3101 = n2742 & ~n2930 ;
  assign n3102 = n2830 & n3101 ;
  assign n3108 = n3107 ^ n3102 ;
  assign n3109 = n3108 ^ n2742 ;
  assign n3118 = n3117 ^ n3109 ;
  assign n3089 = n2005 & ~n2180 ;
  assign n3090 = n3089 ^ n2739 ;
  assign n3119 = n3118 ^ n3090 ;
  assign n3120 = n3088 & n3119 ;
  assign n3121 = n3120 ^ n3088 ;
  assign n3122 = n3121 ^ n3119 ;
  assign n3168 = n2791 & n2955 ;
  assign n3169 = n3168 ^ n2791 ;
  assign n3166 = n2791 & n2940 ;
  assign n3167 = n3166 ^ n2791 ;
  assign n3170 = n3169 ^ n3167 ;
  assign n3164 = n2791 & ~n2930 ;
  assign n3165 = n2830 & n3164 ;
  assign n3171 = n3170 ^ n3165 ;
  assign n3159 = n2773 & n2955 ;
  assign n3160 = n3159 ^ n2773 ;
  assign n3157 = n2773 & n2940 ;
  assign n3158 = n3157 ^ n2773 ;
  assign n3161 = n3160 ^ n3158 ;
  assign n3155 = n2773 & ~n2930 ;
  assign n3156 = n2830 & n3155 ;
  assign n3162 = n3161 ^ n3156 ;
  assign n3163 = n3162 ^ n2773 ;
  assign n3172 = n3171 ^ n3163 ;
  assign n3123 = n2049 & ~n2180 ;
  assign n3124 = n3123 ^ n2770 ;
  assign n3173 = n3172 ^ n3124 ;
  assign n3187 = n2822 & n2955 ;
  assign n3188 = n3187 ^ n2822 ;
  assign n3185 = n2822 & n2940 ;
  assign n3186 = n3185 ^ n2822 ;
  assign n3189 = n3188 ^ n3186 ;
  assign n3183 = n2822 & ~n2930 ;
  assign n3184 = n2830 & n3183 ;
  assign n3190 = n3189 ^ n3184 ;
  assign n3178 = n2798 & n2955 ;
  assign n3179 = n3178 ^ n2798 ;
  assign n3176 = n2798 & n2940 ;
  assign n3177 = n3176 ^ n2798 ;
  assign n3180 = n3179 ^ n3177 ;
  assign n3174 = n2798 & ~n2930 ;
  assign n3175 = n2830 & n3174 ;
  assign n3181 = n3180 ^ n3175 ;
  assign n3182 = n3181 ^ n2798 ;
  assign n3191 = n3190 ^ n3182 ;
  assign n3128 = n2054 & ~n2180 ;
  assign n3129 = n3128 ^ n2795 ;
  assign n3192 = n3191 ^ n3129 ;
  assign n3193 = n3173 & n3192 ;
  assign n3194 = n3193 ^ n3173 ;
  assign n3195 = n3194 ^ n3192 ;
  assign n3196 = n3122 & n3195 ;
  assign n3197 = n3196 ^ n3122 ;
  assign n3198 = n3197 ^ n3195 ;
  assign n3199 = n3066 & n3198 ;
  assign n3200 = n3199 ^ n3066 ;
  assign n3201 = n3200 ^ n3198 ;
  assign n3021 = n2830 & ~n2930 ;
  assign n3022 = n3021 ^ n2955 ;
  assign n3023 = n3022 ^ n2940 ;
  assign n3145 = ~n2791 & n3124 ;
  assign n3146 = n3023 & n3145 ;
  assign n3134 = ~n2822 & n3129 ;
  assign n3141 = ~n2791 & n3134 ;
  assign n3142 = n3023 & n3141 ;
  assign n3130 = ~n2798 & n3129 ;
  assign n3138 = ~n2773 & n3130 ;
  assign n3139 = n3023 & n3138 ;
  assign n3140 = n3139 ^ n3138 ;
  assign n3143 = n3142 ^ n3140 ;
  assign n3135 = n3124 & n3134 ;
  assign n3136 = n3023 & n3135 ;
  assign n3131 = n3124 & n3130 ;
  assign n3132 = n3023 & n3131 ;
  assign n3133 = n3132 ^ n3131 ;
  assign n3137 = n3136 ^ n3133 ;
  assign n3144 = n3143 ^ n3137 ;
  assign n3147 = n3146 ^ n3144 ;
  assign n3125 = ~n2773 & n3124 ;
  assign n3126 = n3023 & n3125 ;
  assign n3127 = n3126 ^ n3125 ;
  assign n3148 = n3147 ^ n3127 ;
  assign n3149 = n3122 & n3148 ;
  assign n3150 = n3149 ^ n3148 ;
  assign n3094 = n2760 & n3090 ;
  assign n3095 = n3023 & n3094 ;
  assign n3091 = n2742 & n3090 ;
  assign n3092 = n3023 & n3091 ;
  assign n3093 = n3092 ^ n3091 ;
  assign n3096 = n3095 ^ n3093 ;
  assign n3097 = n3096 ^ n3090 ;
  assign n3098 = n3088 & n3097 ;
  assign n3099 = n3098 ^ n3097 ;
  assign n3087 = n3068 & ~n3086 ;
  assign n3100 = n3099 ^ n3087 ;
  assign n3151 = n3150 ^ n3100 ;
  assign n3152 = n3066 & n3151 ;
  assign n3153 = n3152 ^ n3151 ;
  assign n3038 = ~n2988 & n2990 ;
  assign n3039 = ~n2969 & n3038 ;
  assign n3029 = n2923 & n3025 ;
  assign n3030 = n3023 & n3029 ;
  assign n3026 = n2905 & n3025 ;
  assign n3027 = n3023 & n3026 ;
  assign n3028 = n3027 ^ n3026 ;
  assign n3031 = n3030 ^ n3028 ;
  assign n3032 = n3031 ^ n3025 ;
  assign n3033 = n3020 & n3032 ;
  assign n3034 = n3033 ^ n3032 ;
  assign n3019 = n3000 & ~n3018 ;
  assign n3035 = n3034 ^ n3019 ;
  assign n3036 = n2998 & n3035 ;
  assign n3037 = n3036 ^ n3035 ;
  assign n3040 = n3039 ^ n3037 ;
  assign n2991 = n2183 & n2990 ;
  assign n2992 = ~n2988 & n2991 ;
  assign n2970 = n2183 & ~n2969 ;
  assign n2993 = n2992 ^ n2970 ;
  assign n3041 = n3040 ^ n2993 ;
  assign n3154 = n3153 ^ n3041 ;
  assign n3202 = n3201 ^ n3154 ;
  assign n3206 = n2969 & n3202 ;
  assign n3207 = n3206 ^ n2969 ;
  assign n3203 = n2183 & n3202 ;
  assign n3204 = n3203 ^ n2183 ;
  assign n3205 = n3204 ^ n2183 ;
  assign n3208 = n3207 ^ n3205 ;
  assign n3212 = n2988 & n3202 ;
  assign n3213 = n3212 ^ n2988 ;
  assign n3209 = n2990 & n3202 ;
  assign n3210 = n3209 ^ n2990 ;
  assign n3211 = n3210 ^ n2990 ;
  assign n3214 = n3213 ^ n3211 ;
  assign n3218 = n3018 & n3202 ;
  assign n3219 = n3218 ^ n3018 ;
  assign n3215 = n3000 & n3202 ;
  assign n3216 = n3215 ^ n3000 ;
  assign n3217 = n3216 ^ n3000 ;
  assign n3220 = n3219 ^ n3217 ;
  assign n3224 = n3059 & n3202 ;
  assign n3225 = n3224 ^ n3059 ;
  assign n3221 = n3025 & n3202 ;
  assign n3222 = n3221 ^ n3025 ;
  assign n3223 = n3222 ^ n3025 ;
  assign n3226 = n3225 ^ n3223 ;
  assign n3230 = n3086 & n3202 ;
  assign n3231 = n3230 ^ n3086 ;
  assign n3227 = n3068 & n3202 ;
  assign n3228 = n3227 ^ n3068 ;
  assign n3229 = n3228 ^ n3068 ;
  assign n3232 = n3231 ^ n3229 ;
  assign n3236 = n3118 & n3202 ;
  assign n3237 = n3236 ^ n3118 ;
  assign n3233 = n3090 & n3202 ;
  assign n3234 = n3233 ^ n3090 ;
  assign n3235 = n3234 ^ n3090 ;
  assign n3238 = n3237 ^ n3235 ;
  assign n3242 = n3172 & n3202 ;
  assign n3243 = n3242 ^ n3172 ;
  assign n3239 = n3124 & n3202 ;
  assign n3240 = n3239 ^ n3124 ;
  assign n3241 = n3240 ^ n3124 ;
  assign n3244 = n3243 ^ n3241 ;
  assign n3248 = n3191 & n3202 ;
  assign n3249 = n3248 ^ n3191 ;
  assign n3245 = n3129 & n3202 ;
  assign n3246 = n3245 ^ n3129 ;
  assign n3247 = n3246 ^ n3129 ;
  assign n3250 = n3249 ^ n3247 ;
  assign n3251 = n3207 ^ n2969 ;
  assign n3252 = n3251 ^ n3204 ;
  assign n3253 = n3213 ^ n2988 ;
  assign n3254 = n3253 ^ n3210 ;
  assign n3255 = n3219 ^ n3018 ;
  assign n3256 = n3255 ^ n3216 ;
  assign n3257 = n3225 ^ n3059 ;
  assign n3258 = n3257 ^ n3222 ;
  assign n3259 = n3231 ^ n3086 ;
  assign n3260 = n3259 ^ n3228 ;
  assign n3261 = n3237 ^ n3118 ;
  assign n3262 = n3261 ^ n3234 ;
  assign n3263 = n3243 ^ n3172 ;
  assign n3264 = n3263 ^ n3240 ;
  assign n3265 = n3249 ^ n3191 ;
  assign n3266 = n3265 ^ n3246 ;
  assign n3267 = n2851 & ~n3023 ;
  assign n3268 = n3267 ^ n2959 ;
  assign n3269 = n2874 & ~n3023 ;
  assign n3270 = n3269 ^ n2978 ;
  assign n3271 = n2900 & ~n3023 ;
  assign n3272 = n3271 ^ n3008 ;
  assign n3273 = n2923 & ~n3023 ;
  assign n3274 = n3273 ^ n3049 ;
  assign n3275 = n2736 & ~n3023 ;
  assign n3276 = n3275 ^ n3076 ;
  assign n3277 = n2760 & ~n3023 ;
  assign n3278 = n3277 ^ n3108 ;
  assign n3279 = n2791 & ~n3023 ;
  assign n3280 = n3279 ^ n3162 ;
  assign n3281 = n2822 & ~n3023 ;
  assign n3282 = n3281 ^ n3181 ;
  assign n3283 = n2556 & ~n2697 ;
  assign n3284 = n3283 ^ n2722 ;
  assign n3285 = n3284 ^ n2707 ;
  assign n3286 = n2588 & ~n3285 ;
  assign n3287 = n3286 ^ n2841 ;
  assign n3288 = n2621 & ~n3285 ;
  assign n3289 = n3288 ^ n2864 ;
  assign n3290 = n2657 & ~n3285 ;
  assign n3291 = n3290 ^ n2890 ;
  assign n3292 = n2690 & ~n3285 ;
  assign n3293 = n3292 ^ n2913 ;
  assign n3294 = n2441 & ~n3285 ;
  assign n3295 = n3294 ^ n2726 ;
  assign n3296 = n2475 & ~n3285 ;
  assign n3297 = n3296 ^ n2750 ;
  assign n3298 = n2514 & ~n3285 ;
  assign n3299 = n3298 ^ n2781 ;
  assign n3300 = n2548 & ~n3285 ;
  assign n3301 = n3300 ^ n2809 ;
  assign n3303 = n2371 & n2422 ;
  assign n3304 = n3303 ^ n2422 ;
  assign n3305 = n3304 ^ n2415 ;
  assign n3302 = n2350 & ~n2395 ;
  assign n3306 = n3305 ^ n3302 ;
  assign n3307 = n3306 ^ n2408 ;
  assign n3309 = n2352 & ~n3307 ;
  assign n3308 = n2358 & n3307 ;
  assign n3310 = n3309 ^ n3308 ;
  assign n3312 = n2361 & ~n3307 ;
  assign n3311 = n2367 & n3307 ;
  assign n3313 = n3312 ^ n3311 ;
  assign n3315 = n2373 & ~n3307 ;
  assign n3314 = n2379 & n3307 ;
  assign n3316 = n3315 ^ n3314 ;
  assign n3318 = n2382 & ~n3307 ;
  assign n3317 = n2388 & n3307 ;
  assign n3319 = n3318 ^ n3317 ;
  assign n3321 = n2195 & ~n3307 ;
  assign n3320 = n2304 & n3307 ;
  assign n3322 = n3321 ^ n3320 ;
  assign n3324 = n2308 & ~n3307 ;
  assign n3323 = n2314 & n3307 ;
  assign n3325 = n3324 ^ n3323 ;
  assign n3327 = n2325 & ~n3307 ;
  assign n3326 = n2331 & n3307 ;
  assign n3328 = n3327 ^ n3326 ;
  assign n3329 = n2342 & n3307 ;
  assign n3330 = n3329 ^ n2534 ;
  assign n3331 = n2356 ^ n2354 ;
  assign n3332 = n2365 ^ n2363 ;
  assign n3333 = n2377 ^ n2375 ;
  assign n3334 = n2386 ^ n2384 ;
  assign n3335 = n2302 ^ n2300 ;
  assign n3336 = n2312 ^ n2310 ;
  assign n3337 = n2329 ^ n2327 ;
  assign n3338 = n2340 ^ n2338 ;
  assign y0 = n3208 ;
  assign y1 = n3214 ;
  assign y2 = n3220 ;
  assign y3 = n3226 ;
  assign y4 = n3232 ;
  assign y5 = n3238 ;
  assign y6 = n3244 ;
  assign y7 = n3250 ;
  assign y8 = n3252 ;
  assign y9 = n3254 ;
  assign y10 = n3256 ;
  assign y11 = n3258 ;
  assign y12 = n3260 ;
  assign y13 = n3262 ;
  assign y14 = n3264 ;
  assign y15 = n3266 ;
  assign y16 = n3268 ;
  assign y17 = n3270 ;
  assign y18 = n3272 ;
  assign y19 = n3274 ;
  assign y20 = n3276 ;
  assign y21 = n3278 ;
  assign y22 = n3280 ;
  assign y23 = n3282 ;
  assign y24 = n3287 ;
  assign y25 = n3289 ;
  assign y26 = n3291 ;
  assign y27 = n3293 ;
  assign y28 = n3295 ;
  assign y29 = n3297 ;
  assign y30 = n3299 ;
  assign y31 = n3301 ;
  assign y32 = n3310 ;
  assign y33 = n3313 ;
  assign y34 = n3316 ;
  assign y35 = n3319 ;
  assign y36 = n3322 ;
  assign y37 = n3325 ;
  assign y38 = n3328 ;
  assign y39 = n3330 ;
  assign y40 = n3331 ;
  assign y41 = n3332 ;
  assign y42 = n3333 ;
  assign y43 = n3334 ;
  assign y44 = n3335 ;
  assign y45 = n3336 ;
  assign y46 = n3337 ;
  assign y47 = n3338 ;
endmodule
