module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 ;
  assign n8 = x0 & x1 ;
  assign n9 = n8 ^ x0 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = x3 & x4 ;
  assign n12 = ~n10 & n11 ;
  assign n13 = n12 ^ n11 ;
  assign n19 = x2 & x3 ;
  assign n20 = x4 & n19 ;
  assign n14 = n11 ^ x3 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = x1 & x2 ;
  assign n17 = n15 & n16 ;
  assign n18 = n17 ^ n16 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n13 & n21 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = n23 ^ n21 ;
  assign n53 = x4 ^ x2 ;
  assign n59 = ~x1 & ~n53 ;
  assign n61 = x4 ^ x0 ;
  assign n62 = n61 ^ x4 ;
  assign n26 = x4 ^ x3 ;
  assign n60 = n26 ^ x4 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n62 ^ x4 ;
  assign n65 = n63 & ~n64 ;
  assign n66 = n65 ^ n62 ;
  assign n67 = n59 & ~n66 ;
  assign n25 = x3 ^ x1 ;
  assign n29 = n25 ^ x4 ;
  assign n30 = x1 & n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n31 ^ x0 ;
  assign n46 = n25 ^ x2 ;
  assign n44 = n31 ^ x3 ;
  assign n45 = n44 ^ x4 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n32 & n47 ;
  assign n49 = n48 ^ n47 ;
  assign n33 = n32 ^ x4 ;
  assign n28 = x2 ^ x1 ;
  assign n34 = n33 ^ n28 ;
  assign n40 = x3 & n34 ;
  assign n41 = n40 ^ x3 ;
  assign n38 = n31 & n34 ;
  assign n39 = n38 ^ n31 ;
  assign n42 = n41 ^ n39 ;
  assign n35 = x0 & n34 ;
  assign n36 = n35 ^ x0 ;
  assign n37 = n36 ^ n34 ;
  assign n43 = n42 ^ n37 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n50 ^ n31 ;
  assign n52 = n51 ^ x1 ;
  assign n54 = n53 ^ n52 ;
  assign n57 = n49 & ~n54 ;
  assign n58 = n57 ^ n54 ;
  assign n68 = n67 ^ n58 ;
  assign n55 = x0 & ~n54 ;
  assign n56 = n55 ^ n54 ;
  assign n69 = n68 ^ n56 ;
  assign n70 = n69 ^ n43 ;
  assign n71 = n70 ^ n49 ;
  assign n72 = n71 ^ n30 ;
  assign n73 = n72 ^ n53 ;
  assign n27 = n26 ^ n25 ;
  assign n74 = n73 ^ n27 ;
  assign n82 = n16 ^ x1 ;
  assign n83 = n14 & n82 ;
  assign n77 = n11 ^ x4 ;
  assign n78 = x0 & x2 ;
  assign n79 = n78 ^ x0 ;
  assign n80 = n79 ^ x2 ;
  assign n81 = n77 & ~n80 ;
  assign n84 = n83 ^ n81 ;
  assign n75 = ~x2 & x4 ;
  assign n76 = ~n10 & n75 ;
  assign n85 = n84 ^ n76 ;
  assign n86 = n82 ^ x2 ;
  assign n87 = n86 ^ x4 ;
  assign n88 = x3 & n87 ;
  assign n89 = n88 ^ x3 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n90 ^ n86 ;
  assign n92 = x0 & n11 ;
  assign n93 = n91 & n92 ;
  assign n94 = n93 ^ n91 ;
  assign n97 = x5 ^ x0 ;
  assign n98 = n97 ^ x4 ;
  assign n99 = n98 ^ x5 ;
  assign n100 = n99 ^ x4 ;
  assign n101 = n100 ^ x5 ;
  assign n102 = n101 ^ x4 ;
  assign n148 = x6 & n99 ;
  assign n149 = n148 ^ x6 ;
  assign n150 = n149 ^ n99 ;
  assign n151 = n102 & ~n150 ;
  assign n103 = n102 ^ x3 ;
  assign n106 = x4 & n103 ;
  assign n107 = n106 ^ n103 ;
  assign n104 = x6 & n103 ;
  assign n105 = n104 ^ n103 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n108 ^ x4 ;
  assign n110 = n109 ^ x6 ;
  assign n111 = n110 ^ n103 ;
  assign n145 = n99 & n102 ;
  assign n146 = n145 ^ n102 ;
  assign n147 = n111 & n146 ;
  assign n152 = n151 ^ n147 ;
  assign n144 = x5 & ~n99 ;
  assign n153 = n152 ^ n144 ;
  assign n112 = n111 ^ x6 ;
  assign n113 = n112 ^ n102 ;
  assign n114 = n102 & n113 ;
  assign n115 = n114 ^ n102 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n117 ^ x6 ;
  assign n119 = n118 ^ x5 ;
  assign n154 = n153 ^ n119 ;
  assign n164 = n86 & n154 ;
  assign n165 = n164 ^ n86 ;
  assign n128 = x5 & n111 ;
  assign n139 = n128 ^ x6 ;
  assign n134 = x5 & x6 ;
  assign n135 = n134 ^ x6 ;
  assign n136 = n102 & n135 ;
  assign n137 = n136 ^ n135 ;
  assign n130 = x5 & n102 ;
  assign n131 = n130 ^ n102 ;
  assign n132 = n111 & n131 ;
  assign n133 = n132 ^ n131 ;
  assign n138 = n137 ^ n133 ;
  assign n140 = n139 ^ n138 ;
  assign n126 = x6 & n102 ;
  assign n127 = n111 & n126 ;
  assign n129 = n128 ^ n127 ;
  assign n141 = n140 ^ n129 ;
  assign n162 = n86 & n141 ;
  assign n163 = n162 ^ n86 ;
  assign n166 = n165 ^ n163 ;
  assign n120 = n101 ^ x6 ;
  assign n121 = n120 ^ n26 ;
  assign n122 = n99 & n121 ;
  assign n123 = n122 ^ n99 ;
  assign n160 = n86 & n123 ;
  assign n161 = n119 & n160 ;
  assign n167 = n166 ^ n161 ;
  assign n155 = x2 & n154 ;
  assign n156 = n155 ^ x2 ;
  assign n142 = x2 & n141 ;
  assign n143 = n142 ^ x2 ;
  assign n157 = n156 ^ n143 ;
  assign n124 = x2 & n123 ;
  assign n125 = n119 & n124 ;
  assign n158 = n157 ^ n125 ;
  assign n159 = n158 ^ x2 ;
  assign n168 = n167 ^ n159 ;
  assign n95 = n77 & n78 ;
  assign n96 = n95 ^ x2 ;
  assign n169 = n168 ^ n96 ;
  assign n170 = n16 & n77 ;
  assign n171 = n170 ^ n16 ;
  assign n172 = n171 ^ x1 ;
  assign n173 = n19 ^ x3 ;
  assign n174 = x4 & x6 ;
  assign n175 = n174 ^ x4 ;
  assign n176 = n173 & n175 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = n172 & n177 ;
  assign n179 = n178 ^ n82 ;
  assign n180 = n179 ^ n172 ;
  assign n183 = n26 & n53 ;
  assign n184 = n183 ^ n26 ;
  assign n185 = n184 ^ x4 ;
  assign n186 = n185 ^ x2 ;
  assign n187 = n185 & n186 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = n188 ^ n185 ;
  assign n182 = n8 & n11 ;
  assign n190 = n189 ^ n182 ;
  assign n191 = n190 ^ n11 ;
  assign n192 = x2 & n191 ;
  assign n193 = n192 ^ x2 ;
  assign n194 = n193 ^ n191 ;
  assign n181 = ~n8 & n11 ;
  assign n195 = n194 ^ n181 ;
  assign n196 = n195 ^ n188 ;
  assign n197 = n196 ^ n182 ;
  assign n198 = n197 ^ n11 ;
  assign n208 = x0 & x3 ;
  assign n209 = n208 ^ x3 ;
  assign n210 = x4 & n209 ;
  assign n211 = n210 ^ x4 ;
  assign n212 = n211 ^ x4 ;
  assign n213 = n86 & n212 ;
  assign n214 = n213 ^ n212 ;
  assign n200 = x1 ^ x0 ;
  assign n201 = n200 ^ x1 ;
  assign n199 = x4 ^ x1 ;
  assign n202 = n201 ^ n199 ;
  assign n203 = n199 ^ x1 ;
  assign n204 = n202 & n203 ;
  assign n205 = n204 ^ n199 ;
  assign n206 = x2 & ~n26 ;
  assign n207 = n205 & n206 ;
  assign n215 = n214 ^ n207 ;
  assign n221 = x0 & n77 ;
  assign n222 = n221 ^ n77 ;
  assign n223 = n82 & n222 ;
  assign n224 = n223 ^ n82 ;
  assign n217 = x2 & x4 ;
  assign n218 = n217 ^ x2 ;
  assign n216 = n19 ^ x2 ;
  assign n219 = n218 ^ n216 ;
  assign n220 = x1 & ~n219 ;
  assign n225 = n224 ^ n220 ;
  assign n227 = n11 & ~n86 ;
  assign n228 = n227 ^ n223 ;
  assign n226 = ~n15 & n16 ;
  assign n229 = n228 ^ n226 ;
  assign n233 = n8 ^ x1 ;
  assign n234 = n77 & n233 ;
  assign n235 = n234 ^ n77 ;
  assign n236 = x2 & n235 ;
  assign n237 = n236 ^ n235 ;
  assign n231 = ~x1 & x4 ;
  assign n232 = n173 & ~n231 ;
  assign n238 = n237 ^ n232 ;
  assign n230 = x2 & n77 ;
  assign n239 = n238 ^ n230 ;
  assign n240 = x0 & n15 ;
  assign n241 = n240 ^ x0 ;
  assign n242 = n241 ^ n15 ;
  assign n243 = n86 & ~n242 ;
  assign n244 = n243 ^ n242 ;
  assign n251 = x1 & x3 ;
  assign n252 = n251 ^ x1 ;
  assign n253 = x2 & ~x4 ;
  assign n254 = ~n252 & n253 ;
  assign n245 = ~n10 & n77 ;
  assign n246 = n245 ^ n77 ;
  assign n247 = n246 ^ x3 ;
  assign n248 = x2 & n247 ;
  assign n249 = n248 ^ x2 ;
  assign n250 = n249 ^ n247 ;
  assign n255 = n254 ^ n250 ;
  assign n256 = ~n15 & n78 ;
  assign n257 = ~x0 & x2 ;
  assign n258 = ~n15 & n257 ;
  assign n259 = x1 & n14 ;
  assign n260 = n259 ^ n14 ;
  assign n261 = n257 & n260 ;
  assign n262 = n261 ^ n257 ;
  assign n263 = n262 ^ n257 ;
  assign n264 = n9 & n14 ;
  assign n265 = x2 & n264 ;
  assign n266 = x2 & n14 ;
  assign n267 = n8 & n266 ;
  assign n268 = n233 & n266 ;
  assign n269 = x2 & n15 ;
  assign n270 = n269 ^ x2 ;
  assign n280 = x2 & n182 ;
  assign n279 = x2 & ~n11 ;
  assign n281 = n280 ^ n279 ;
  assign n273 = n8 & n173 ;
  assign n274 = x4 & x5 ;
  assign n275 = n274 ^ x4 ;
  assign n276 = n273 & n275 ;
  assign n277 = n276 ^ n273 ;
  assign n271 = n265 ^ x2 ;
  assign n272 = n271 ^ n264 ;
  assign n278 = n277 ^ n272 ;
  assign n282 = n281 ^ n278 ;
  assign n288 = ~x1 & x3 ;
  assign n289 = x4 & n79 ;
  assign n290 = n289 ^ n79 ;
  assign n291 = n288 & n290 ;
  assign n283 = n11 & n79 ;
  assign n284 = x1 & x5 ;
  assign n285 = x6 & n284 ;
  assign n286 = n285 ^ n284 ;
  assign n287 = n283 & n286 ;
  assign n292 = n291 ^ n287 ;
  assign n302 = n280 ^ x2 ;
  assign n303 = n302 ^ n279 ;
  assign n293 = n11 & n134 ;
  assign n294 = n293 ^ n11 ;
  assign n295 = n294 ^ x3 ;
  assign n298 = x2 & n8 ;
  assign n299 = n295 & n298 ;
  assign n300 = n299 ^ n295 ;
  assign n296 = n8 & n295 ;
  assign n297 = n296 ^ n295 ;
  assign n301 = n300 ^ n297 ;
  assign n304 = n303 ^ n301 ;
  assign n305 = n77 ^ x2 ;
  assign n306 = n200 ^ x2 ;
  assign n307 = n200 & n306 ;
  assign n308 = n307 ^ x2 ;
  assign n309 = ~n305 & n308 ;
  assign n310 = n309 ^ n307 ;
  assign n311 = n310 ^ n77 ;
  assign n312 = x1 & n77 ;
  assign n313 = n312 ^ n77 ;
  assign n314 = n79 & n313 ;
  assign y0 = n24 ;
  assign y1 = ~n74 ;
  assign y2 = n85 ;
  assign y3 = n94 ;
  assign y4 = n169 ;
  assign y5 = n180 ;
  assign y6 = n198 ;
  assign y7 = n215 ;
  assign y8 = n225 ;
  assign y9 = n229 ;
  assign y10 = n239 ;
  assign y11 = ~n244 ;
  assign y12 = n255 ;
  assign y13 = n256 ;
  assign y14 = n258 ;
  assign y15 = n263 ;
  assign y16 = n265 ;
  assign y17 = n267 ;
  assign y18 = n268 ;
  assign y19 = n270 ;
  assign y20 = n282 ;
  assign y21 = n292 ;
  assign y22 = n304 ;
  assign y23 = ~1'b0 ;
  assign y24 = n311 ;
  assign y25 = n314 ;
endmodule
