module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 ;
  assign n33 = ~x0 & ~x1 ;
  assign n34 = x2 & x3 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = x4 & x5 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n36 & n39 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n33 & n42 ;
  assign n44 = n43 ^ n33 ;
  assign n45 = x10 & x11 ;
  assign n46 = n45 ^ x10 ;
  assign n47 = n46 ^ x11 ;
  assign n48 = x13 & x14 ;
  assign n49 = n48 ^ x13 ;
  assign n50 = n49 ^ x14 ;
  assign n51 = n47 & n50 ;
  assign n52 = n51 ^ n47 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = x6 & x7 ;
  assign n55 = n54 ^ x6 ;
  assign n56 = n55 ^ x7 ;
  assign n57 = x8 & x9 ;
  assign n58 = n57 ^ x8 ;
  assign n59 = n58 ^ x9 ;
  assign n60 = n56 & n59 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n53 & n62 ;
  assign n64 = n63 ^ n53 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n44 & ~n65 ;
  assign n67 = x21 & x22 ;
  assign n68 = n67 ^ x21 ;
  assign n69 = n68 ^ x22 ;
  assign n70 = x20 & x23 ;
  assign n71 = n70 ^ x20 ;
  assign n72 = n71 ^ x23 ;
  assign n73 = n69 & ~n72 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~x24 & ~x25 ;
  assign n76 = ~n74 & n75 ;
  assign n77 = x16 & x17 ;
  assign n78 = n77 ^ x16 ;
  assign n79 = n78 ^ x17 ;
  assign n80 = x18 & n79 ;
  assign n81 = n80 ^ x18 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = x12 & x15 ;
  assign n84 = n83 ^ x12 ;
  assign n85 = n84 ^ x15 ;
  assign n86 = x19 & ~n85 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n82 & ~n87 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ n76 ;
  assign n91 = n76 & ~n90 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n93 ^ n66 ;
  assign n95 = n66 & n94 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = n96 ^ n92 ;
  assign n98 = n97 ^ n89 ;
  assign n99 = ~x28 & ~x29 ;
  assign n100 = ~x30 & ~x31 ;
  assign n101 = n99 & n100 ;
  assign n104 = x26 & ~x27 ;
  assign n105 = n101 & n104 ;
  assign n102 = ~x26 & ~x27 ;
  assign n103 = n101 & n102 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = n98 & n106 ;
  assign n108 = n107 ^ n103 ;
  assign n109 = ~n82 & ~n85 ;
  assign n110 = n66 & n109 ;
  assign n111 = ~x19 & ~n74 ;
  assign n112 = x24 & ~x25 ;
  assign n113 = n112 ^ n75 ;
  assign n114 = n111 & n113 ;
  assign n115 = n110 & n114 ;
  assign n116 = n115 ^ n75 ;
  assign n117 = n108 & n116 ;
  assign n118 = n117 ^ n108 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = n119 ^ n108 ;
  assign n121 = n120 ^ n116 ;
  assign n122 = ~x16 & ~x17 ;
  assign n123 = x18 & ~n85 ;
  assign n124 = n122 & n123 ;
  assign n125 = n66 & n124 ;
  assign n126 = n125 ^ x18 ;
  assign n127 = n111 ^ n109 ;
  assign n128 = ~n111 & ~n127 ;
  assign n129 = n128 ^ n111 ;
  assign n130 = n129 ^ n66 ;
  assign n131 = n109 ^ n66 ;
  assign n132 = ~n130 & n131 ;
  assign n133 = n132 ^ n128 ;
  assign n134 = n133 ^ n66 ;
  assign n135 = n126 & ~n134 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = ~n121 & ~n136 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n33 & ~n85 ;
  assign n140 = ~n42 & n139 ;
  assign n141 = ~n65 & n140 ;
  assign n142 = n141 ^ x16 ;
  assign n143 = ~x17 & ~n142 ;
  assign n144 = ~n138 & n143 ;
  assign n145 = n142 ^ n136 ;
  assign n146 = ~n142 & ~n145 ;
  assign n147 = n146 ^ n136 ;
  assign n148 = n147 ^ n121 ;
  assign n149 = ~n121 & ~n148 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = n150 ^ n136 ;
  assign n152 = n151 ^ n138 ;
  assign n153 = x17 & n152 ;
  assign n154 = n98 & n103 ;
  assign n155 = n154 ^ n103 ;
  assign n156 = x24 & ~n74 ;
  assign n157 = n156 ^ n74 ;
  assign n158 = n157 ^ n89 ;
  assign n159 = ~n157 & n158 ;
  assign n160 = n159 ^ n158 ;
  assign n161 = n160 ^ n89 ;
  assign n162 = n161 ^ n66 ;
  assign n163 = n66 & ~n162 ;
  assign n164 = n163 ^ n162 ;
  assign n165 = n164 ^ n160 ;
  assign n166 = n165 ^ n89 ;
  assign n167 = x25 & n166 ;
  assign n168 = n167 ^ x25 ;
  assign n169 = n155 & n168 ;
  assign n170 = n169 ^ n155 ;
  assign n171 = x19 & ~n110 ;
  assign n172 = n66 & ~n89 ;
  assign n173 = ~n157 & ~n172 ;
  assign n174 = ~n171 & n173 ;
  assign n175 = n170 & n174 ;
  assign n176 = x16 & n141 ;
  assign n177 = n176 ^ n141 ;
  assign n178 = x17 & ~n177 ;
  assign n179 = n122 & n141 ;
  assign n180 = ~x18 & ~n179 ;
  assign n181 = ~n178 & n180 ;
  assign n182 = n175 & n181 ;
  assign n183 = n153 & n182 ;
  assign n184 = n183 ^ n153 ;
  assign n185 = n184 ^ n152 ;
  assign n186 = n185 ^ n182 ;
  assign n187 = n182 ^ n138 ;
  assign n188 = ~n144 & ~n187 ;
  assign n189 = ~n138 & n175 ;
  assign n190 = n181 ^ n138 ;
  assign n191 = n175 & ~n190 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = n192 ^ n175 ;
  assign n194 = n193 ^ n181 ;
  assign n195 = n189 & ~n194 ;
  assign n196 = n195 ^ n194 ;
  assign n197 = ~n138 & ~n175 ;
  assign n198 = x23 & ~n69 ;
  assign n199 = n198 ^ n69 ;
  assign n200 = n172 ^ x20 ;
  assign n201 = n199 & n200 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = ~n121 & ~n203 ;
  assign n205 = n204 ^ n203 ;
  assign n206 = n197 & ~n205 ;
  assign n207 = n206 ^ n175 ;
  assign n208 = n207 ^ n205 ;
  assign n209 = n175 & n205 ;
  assign n210 = ~x22 & ~x23 ;
  assign n211 = ~x24 & n210 ;
  assign n212 = n66 ^ x20 ;
  assign n213 = n89 ^ x20 ;
  assign n214 = n89 & n213 ;
  assign n215 = n214 ^ x20 ;
  assign n216 = ~n212 & n215 ;
  assign n217 = n216 ^ n214 ;
  assign n218 = n217 ^ n66 ;
  assign n219 = n218 ^ x21 ;
  assign n220 = n219 ^ n211 ;
  assign n221 = ~n211 & ~n220 ;
  assign n222 = n221 ^ n219 ;
  assign n223 = n222 ^ n170 ;
  assign n224 = ~n170 & ~n223 ;
  assign n225 = n224 ^ n221 ;
  assign n226 = n225 ^ n219 ;
  assign n227 = n209 & ~n226 ;
  assign n228 = n227 ^ n205 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = n170 ^ n116 ;
  assign n231 = ~x24 & ~n219 ;
  assign n232 = n231 ^ n116 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = n233 ^ n116 ;
  assign n235 = ~n230 & n234 ;
  assign n236 = n235 ^ n233 ;
  assign n237 = n236 ^ n170 ;
  assign n238 = n237 ^ n231 ;
  assign n239 = n205 & n238 ;
  assign n240 = n239 ^ n238 ;
  assign n241 = n240 ^ n205 ;
  assign n242 = n241 ^ n238 ;
  assign n243 = ~n121 & ~n231 ;
  assign n244 = x21 & n218 ;
  assign n245 = n244 ^ n218 ;
  assign n246 = n245 ^ x22 ;
  assign n247 = x23 & n246 ;
  assign n248 = n247 ^ n246 ;
  assign n249 = n248 ^ x23 ;
  assign n250 = n243 & ~n249 ;
  assign n251 = n250 ^ n249 ;
  assign n252 = n242 & n251 ;
  assign n253 = n252 ^ n242 ;
  assign n254 = ~x22 & n245 ;
  assign n255 = x23 & ~n254 ;
  assign n256 = n110 & n111 ;
  assign n257 = ~x24 & ~n256 ;
  assign n258 = n170 & n257 ;
  assign n259 = ~n255 & n258 ;
  assign n260 = n249 & n259 ;
  assign n261 = n121 & ~n259 ;
  assign n262 = n116 & n170 ;
  assign n263 = n262 ^ n170 ;
  assign n264 = n108 & ~n116 ;
  assign n265 = ~n170 & n264 ;
  assign n266 = x26 & n98 ;
  assign n267 = n266 ^ n98 ;
  assign n268 = ~n104 & ~n267 ;
  assign n269 = ~x27 & n98 ;
  assign n270 = n101 & ~n269 ;
  assign n271 = ~n268 & n270 ;
  assign n272 = x27 & ~x28 ;
  assign n273 = ~n267 & n272 ;
  assign n274 = n98 & n102 ;
  assign n275 = x28 & n274 ;
  assign n276 = ~n273 & ~n275 ;
  assign n277 = ~x29 & n100 ;
  assign n278 = ~n276 & n277 ;
  assign n279 = x29 & ~n274 ;
  assign n280 = ~n99 & n100 ;
  assign n281 = ~n275 & n280 ;
  assign n282 = ~n279 & n281 ;
  assign n283 = n275 ^ n274 ;
  assign n285 = x29 & n100 ;
  assign n284 = x30 & ~x31 ;
  assign n286 = n285 ^ n284 ;
  assign n288 = n286 ^ x29 ;
  assign n287 = n286 ^ n284 ;
  assign n289 = n288 ^ n287 ;
  assign n290 = n287 ^ n286 ;
  assign n291 = n289 & n290 ;
  assign n292 = n291 ^ n287 ;
  assign n293 = n283 & n292 ;
  assign n294 = n293 ^ n286 ;
  assign n295 = n294 ^ n284 ;
  assign n296 = n99 & n102 ;
  assign n297 = n98 & n296 ;
  assign n298 = n297 ^ x31 ;
  assign n299 = n297 ^ x30 ;
  assign n300 = n298 & n299 ;
  assign n301 = n300 ^ n299 ;
  assign y0 = n144 ;
  assign y1 = n186 ;
  assign y2 = n188 ;
  assign y3 = ~n196 ;
  assign y4 = ~n208 ;
  assign y5 = n229 ;
  assign y6 = n253 ;
  assign y7 = n260 ;
  assign y8 = n261 ;
  assign y9 = n263 ;
  assign y10 = n265 ;
  assign y11 = n271 ;
  assign y12 = n278 ;
  assign y13 = n282 ;
  assign y14 = n295 ;
  assign y15 = n301 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
  assign y30 = 1'b0 ;
  assign y31 = 1'b0 ;
endmodule
