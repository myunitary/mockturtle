module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 ;
  assign n150 = x4 & x19 ;
  assign n151 = n150 ^ x4 ;
  assign n152 = n151 ^ x19 ;
  assign n153 = ~x16 & ~x18 ;
  assign n154 = ~n152 & n153 ;
  assign n148 = ~x5 & ~x22 ;
  assign n155 = ~x6 & ~x12 ;
  assign n156 = ~x17 & n155 ;
  assign n157 = n148 & n156 ;
  assign n158 = n154 & n157 ;
  assign n159 = ~x8 & ~x21 ;
  assign n160 = ~x7 & ~x13 ;
  assign n174 = x14 & n160 ;
  assign n175 = n159 & n174 ;
  assign n168 = ~x8 & ~x13 ;
  assign n169 = ~x21 & n168 ;
  assign n167 = ~x21 & n160 ;
  assign n170 = n169 ^ n167 ;
  assign n163 = ~x7 & ~x8 ;
  assign n165 = x13 & n163 ;
  assign n164 = x21 & n163 ;
  assign n166 = n165 ^ n164 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = ~x10 & ~x14 ;
  assign n173 = n171 & n172 ;
  assign n176 = n175 ^ n173 ;
  assign n161 = x10 & n160 ;
  assign n162 = n159 & n161 ;
  assign n177 = n176 ^ n162 ;
  assign n178 = ~x9 & ~x11 ;
  assign n183 = n177 & n178 ;
  assign n184 = n158 & n183 ;
  assign n179 = ~x56 & n178 ;
  assign n180 = ~n148 & n179 ;
  assign n181 = n177 & n180 ;
  assign n182 = n158 & n181 ;
  assign n185 = n184 ^ n182 ;
  assign n186 = n185 ^ n179 ;
  assign n149 = ~x56 & n148 ;
  assign n187 = n186 ^ n149 ;
  assign n190 = ~x14 & ~x22 ;
  assign n191 = n160 & n190 ;
  assign n192 = n178 & n191 ;
  assign n193 = ~x17 & ~x21 ;
  assign n194 = ~x8 & n193 ;
  assign n195 = ~x5 & n155 ;
  assign n196 = n194 & n195 ;
  assign n197 = n192 & n196 ;
  assign n198 = ~x0 & x54 ;
  assign n199 = n154 & n198 ;
  assign n200 = n197 & n199 ;
  assign n201 = ~n187 & n200 ;
  assign n189 = x0 & ~x54 ;
  assign n202 = n201 ^ n189 ;
  assign n188 = x54 & ~n187 ;
  assign n203 = n202 ^ n188 ;
  assign n204 = ~x3 & ~x129 ;
  assign n205 = ~n203 & n204 ;
  assign n206 = ~x5 & ~x6 ;
  assign n207 = ~x7 & ~x12 ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = ~x13 & ~n208 ;
  assign n210 = ~x5 & ~x7 ;
  assign n211 = n210 ^ n155 ;
  assign n212 = n209 & n211 ;
  assign n213 = x13 & n155 ;
  assign n214 = n210 & n213 ;
  assign n215 = ~x9 & ~n214 ;
  assign n216 = ~n212 & n215 ;
  assign n217 = n160 & n195 ;
  assign n218 = x9 & ~n217 ;
  assign n219 = ~x10 & x54 ;
  assign n220 = n190 & n219 ;
  assign n221 = ~x8 & ~x11 ;
  assign n222 = n193 & n221 ;
  assign n223 = n220 & n222 ;
  assign n224 = n154 & n223 ;
  assign n225 = ~n218 & n224 ;
  assign n226 = ~n216 & n225 ;
  assign n227 = n160 & n206 ;
  assign n228 = n154 & n227 ;
  assign n229 = ~x14 & n159 ;
  assign n230 = ~x11 & ~x12 ;
  assign n231 = ~x10 & ~x22 ;
  assign n232 = n230 & n231 ;
  assign n233 = n229 & n232 ;
  assign n234 = n228 & n233 ;
  assign n235 = ~x17 & x54 ;
  assign n236 = ~x1 & n235 ;
  assign n237 = ~n234 & n236 ;
  assign n238 = n237 ^ x1 ;
  assign n239 = n204 & n238 ;
  assign n240 = ~n226 & n239 ;
  assign n241 = n240 ^ n204 ;
  assign n242 = x38 & x50 ;
  assign n243 = n242 ^ x38 ;
  assign n244 = n243 ^ x50 ;
  assign n245 = ~x40 & ~x46 ;
  assign n246 = ~n244 & n245 ;
  assign n247 = x41 & x43 ;
  assign n248 = n247 ^ x41 ;
  assign n249 = n248 ^ x43 ;
  assign n250 = x42 & x44 ;
  assign n251 = n250 ^ x42 ;
  assign n252 = n251 ^ x44 ;
  assign n253 = ~n249 & ~n252 ;
  assign n254 = n246 & n253 ;
  assign n255 = x47 & x48 ;
  assign n256 = n255 ^ x47 ;
  assign n257 = n256 ^ x48 ;
  assign n258 = n254 & ~n257 ;
  assign n259 = x15 & x20 ;
  assign n260 = n259 ^ x15 ;
  assign n261 = n260 ^ x20 ;
  assign n262 = ~x45 & ~n261 ;
  assign n263 = x24 & x49 ;
  assign n264 = n263 ^ x24 ;
  assign n265 = n264 ^ x49 ;
  assign n266 = x82 & ~n265 ;
  assign n267 = n262 & n266 ;
  assign n268 = x122 & x127 ;
  assign n269 = ~x82 & ~n268 ;
  assign n270 = x2 & ~n269 ;
  assign n271 = n267 & n270 ;
  assign n272 = n258 & n271 ;
  assign n273 = n272 ^ n270 ;
  assign n283 = ~x65 & ~n268 ;
  assign n288 = ~x82 & n283 ;
  assign n289 = ~n273 & n288 ;
  assign n290 = n289 ^ n273 ;
  assign n274 = n262 & ~n265 ;
  assign n275 = ~x41 & ~x46 ;
  assign n276 = ~n244 & n275 ;
  assign n277 = ~x43 & ~x47 ;
  assign n278 = ~x2 & ~x48 ;
  assign n279 = n277 & n278 ;
  assign n280 = n276 & n279 ;
  assign n281 = n274 & n280 ;
  assign n282 = ~x40 & ~n252 ;
  assign n284 = x82 & n283 ;
  assign n285 = n282 & n284 ;
  assign n286 = n281 & n285 ;
  assign n287 = ~n273 & n286 ;
  assign n291 = n290 ^ n287 ;
  assign n292 = ~x129 & n291 ;
  assign n297 = x0 & ~x113 ;
  assign n298 = ~x123 & n297 ;
  assign n299 = ~x61 & ~x118 ;
  assign n304 = ~x129 & ~n299 ;
  assign n305 = ~n298 & n304 ;
  assign n306 = n305 ^ x129 ;
  assign n293 = ~x9 & ~x14 ;
  assign n294 = n231 & n293 ;
  assign n295 = ~x12 & n222 ;
  assign n296 = n294 & n295 ;
  assign n300 = ~x129 & n299 ;
  assign n301 = ~n298 & n300 ;
  assign n302 = n228 & n301 ;
  assign n303 = n296 & n302 ;
  assign n307 = n306 ^ n303 ;
  assign n310 = x18 & ~n152 ;
  assign n311 = n310 ^ n152 ;
  assign n312 = ~x16 & x54 ;
  assign n313 = n193 & n312 ;
  assign n314 = ~n311 & n313 ;
  assign n315 = x10 & ~x22 ;
  assign n316 = n221 & n315 ;
  assign n317 = n314 & n316 ;
  assign n318 = n160 & n293 ;
  assign n319 = n195 & n318 ;
  assign n308 = x4 & ~x54 ;
  assign n320 = n204 & ~n308 ;
  assign n321 = n319 & n320 ;
  assign n322 = n317 & n321 ;
  assign n309 = n204 & n308 ;
  assign n323 = n322 ^ n309 ;
  assign n324 = x5 & ~x54 ;
  assign n325 = ~x13 & n294 ;
  assign n326 = ~x59 & n222 ;
  assign n327 = n325 & n326 ;
  assign n328 = n155 & n210 ;
  assign n329 = n312 & n328 ;
  assign n330 = ~x25 & x28 ;
  assign n331 = ~x29 & n330 ;
  assign n332 = ~n311 & n331 ;
  assign n333 = n329 & n332 ;
  assign n334 = n327 & n333 ;
  assign n335 = ~n324 & ~n334 ;
  assign n336 = n204 & ~n335 ;
  assign n337 = x6 & ~x54 ;
  assign n338 = ~x28 & ~x29 ;
  assign n339 = x25 & n338 ;
  assign n340 = ~n311 & n339 ;
  assign n341 = n329 & n340 ;
  assign n342 = n327 & n341 ;
  assign n343 = ~n337 & ~n342 ;
  assign n344 = n204 & ~n343 ;
  assign n345 = x7 & ~x54 ;
  assign n346 = x8 & n314 ;
  assign n347 = ~x11 & n328 ;
  assign n348 = n325 & n347 ;
  assign n349 = n346 & n348 ;
  assign n350 = ~n345 & ~n349 ;
  assign n351 = n204 & ~n350 ;
  assign n352 = x8 & ~x54 ;
  assign n353 = ~x12 & n294 ;
  assign n354 = n227 & n353 ;
  assign n355 = ~n152 & n312 ;
  assign n356 = ~x17 & ~x18 ;
  assign n357 = n221 & n356 ;
  assign n358 = x21 & n357 ;
  assign n359 = n355 & n358 ;
  assign n360 = n354 & n359 ;
  assign n361 = ~n352 & ~n360 ;
  assign n362 = n204 & ~n361 ;
  assign n363 = x9 & ~x54 ;
  assign n364 = ~x8 & n314 ;
  assign n365 = x11 & n328 ;
  assign n366 = n325 & n365 ;
  assign n367 = n364 & n366 ;
  assign n368 = ~n363 & ~n367 ;
  assign n369 = n204 & ~n368 ;
  assign n370 = x10 & ~x54 ;
  assign n371 = ~x9 & ~x18 ;
  assign n372 = n194 & n371 ;
  assign n373 = n231 & n372 ;
  assign n374 = ~x13 & x14 ;
  assign n375 = n355 & n374 ;
  assign n376 = n347 & n375 ;
  assign n377 = n373 & n376 ;
  assign n378 = ~n370 & ~n377 ;
  assign n379 = n204 & ~n378 ;
  assign n382 = ~x10 & ~x11 ;
  assign n383 = x22 & n382 ;
  assign n380 = x11 & ~x54 ;
  assign n384 = n204 & ~n380 ;
  assign n385 = n383 & n384 ;
  assign n386 = n319 & n385 ;
  assign n387 = n364 & n386 ;
  assign n381 = n204 & n380 ;
  assign n388 = n387 ^ n381 ;
  assign n389 = x12 & ~x54 ;
  assign n390 = x18 & n227 ;
  assign n391 = n294 & n355 ;
  assign n392 = n390 & n391 ;
  assign n393 = n295 & n392 ;
  assign n394 = ~n389 & ~n393 ;
  assign n395 = n204 & ~n394 ;
  assign n396 = ~x25 & ~x28 ;
  assign n397 = x29 & n396 ;
  assign n398 = ~x59 & n231 ;
  assign n399 = n397 & n398 ;
  assign n400 = n314 & n399 ;
  assign n401 = x13 & ~x54 ;
  assign n402 = n221 & ~n401 ;
  assign n403 = n319 & n402 ;
  assign n404 = n400 & n403 ;
  assign n405 = n404 ^ n401 ;
  assign n406 = n204 & n405 ;
  assign n407 = x14 & ~x54 ;
  assign n408 = x13 & ~x16 ;
  assign n409 = ~n152 & n408 ;
  assign n410 = n220 & n409 ;
  assign n411 = n347 & n410 ;
  assign n412 = n372 & n411 ;
  assign n413 = ~n407 & ~n412 ;
  assign n414 = n204 & ~n413 ;
  assign n431 = ~n257 & ~n265 ;
  assign n432 = ~x15 & ~x45 ;
  assign n433 = ~n249 & n432 ;
  assign n434 = n431 & n433 ;
  assign n435 = x82 & ~n252 ;
  assign n436 = n246 & n435 ;
  assign n437 = n434 & n436 ;
  assign n438 = n437 ^ x82 ;
  assign n439 = ~x82 & n268 ;
  assign n440 = x15 & n439 ;
  assign n441 = ~x70 & ~n268 ;
  assign n442 = ~n440 & n441 ;
  assign n443 = ~n438 & n442 ;
  assign n444 = n443 ^ n440 ;
  assign n448 = ~x129 & n444 ;
  assign n415 = n276 & n282 ;
  assign n416 = x45 & ~n265 ;
  assign n417 = n416 ^ n265 ;
  assign n418 = ~x48 & n277 ;
  assign n419 = ~n417 & n418 ;
  assign n420 = n415 & n419 ;
  assign n421 = x15 & ~n420 ;
  assign n422 = x15 & ~n265 ;
  assign n423 = n422 ^ n265 ;
  assign n424 = x45 & ~n257 ;
  assign n425 = n424 ^ n257 ;
  assign n426 = ~x2 & ~x20 ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = ~n423 & n427 ;
  assign n429 = n254 & n428 ;
  assign n430 = ~n421 & ~n429 ;
  assign n445 = x82 & ~x129 ;
  assign n446 = ~n444 & n445 ;
  assign n447 = ~n430 & n446 ;
  assign n449 = n448 ^ n447 ;
  assign n450 = x16 & ~x54 ;
  assign n451 = n221 & n314 ;
  assign n452 = x6 & ~x13 ;
  assign n453 = n210 & n452 ;
  assign n454 = n353 & n453 ;
  assign n455 = n451 & n454 ;
  assign n456 = ~n450 & ~n455 ;
  assign n457 = n204 & ~n456 ;
  assign n458 = x17 & ~x54 ;
  assign n459 = ~x25 & x59 ;
  assign n460 = n159 & n459 ;
  assign n461 = n235 & n338 ;
  assign n462 = n460 & n461 ;
  assign n463 = n154 & n462 ;
  assign n464 = n348 & n463 ;
  assign n465 = ~n458 & ~n464 ;
  assign n466 = n204 & ~n465 ;
  assign n469 = n227 & ~n311 ;
  assign n470 = n353 & n469 ;
  assign n471 = x16 & x54 ;
  assign n472 = n222 & n471 ;
  assign n467 = x18 & ~x54 ;
  assign n473 = n204 & ~n467 ;
  assign n474 = n472 & n473 ;
  assign n475 = n470 & n474 ;
  assign n468 = n204 & n467 ;
  assign n476 = n475 ^ n468 ;
  assign n479 = x17 & ~x21 ;
  assign n480 = n221 & n479 ;
  assign n481 = n312 & n480 ;
  assign n477 = x19 & ~x54 ;
  assign n482 = n204 & ~n477 ;
  assign n483 = n481 & n482 ;
  assign n484 = n470 & n483 ;
  assign n478 = n204 & n477 ;
  assign n485 = n484 ^ n478 ;
  assign n487 = ~x46 & ~x50 ;
  assign n488 = x38 & x40 ;
  assign n489 = n488 ^ x38 ;
  assign n490 = n489 ^ x40 ;
  assign n491 = ~n252 & ~n490 ;
  assign n492 = n487 & n491 ;
  assign n493 = ~n249 & ~n265 ;
  assign n494 = ~n425 & n493 ;
  assign n495 = n492 & n494 ;
  assign n498 = ~x2 & ~x15 ;
  assign n499 = ~x20 & x82 ;
  assign n500 = n498 & n499 ;
  assign n501 = n495 & n500 ;
  assign n496 = ~x15 & x82 ;
  assign n497 = n495 & n496 ;
  assign n502 = n501 ^ n497 ;
  assign n486 = x20 & x82 ;
  assign n503 = n502 ^ n486 ;
  assign n504 = x20 & n439 ;
  assign n505 = ~x71 & ~n268 ;
  assign n510 = ~x82 & n505 ;
  assign n511 = ~n504 & n510 ;
  assign n512 = n511 ^ n504 ;
  assign n506 = x82 & ~n261 ;
  assign n507 = n505 & n506 ;
  assign n508 = ~n504 & n507 ;
  assign n509 = n495 & n508 ;
  assign n513 = n512 ^ n509 ;
  assign n514 = ~n503 & ~n513 ;
  assign n515 = ~x129 & ~n514 ;
  assign n516 = x21 & ~x54 ;
  assign n517 = ~x4 & x19 ;
  assign n518 = ~x21 & n517 ;
  assign n519 = n312 & n518 ;
  assign n520 = n357 & n519 ;
  assign n521 = n354 & n520 ;
  assign n522 = ~n516 & ~n521 ;
  assign n523 = n204 & ~n522 ;
  assign n524 = x22 & ~x54 ;
  assign n525 = x5 & ~x6 ;
  assign n526 = ~x14 & n525 ;
  assign n527 = n160 & n230 ;
  assign n528 = n526 & n527 ;
  assign n529 = n355 & n528 ;
  assign n530 = n373 & n529 ;
  assign n531 = ~n524 & ~n530 ;
  assign n532 = n204 & ~n531 ;
  assign n533 = ~x23 & x55 ;
  assign n534 = x61 & ~x129 ;
  assign n535 = ~n533 & n534 ;
  assign n542 = x2 & ~n261 ;
  assign n543 = n542 ^ n261 ;
  assign n553 = ~x49 & ~n543 ;
  assign n554 = x82 & ~n553 ;
  assign n555 = n268 & ~n554 ;
  assign n536 = ~n249 & ~n425 ;
  assign n556 = n246 & ~n252 ;
  assign n557 = n536 & n556 ;
  assign n558 = x82 & ~n557 ;
  assign n559 = ~n555 & ~n558 ;
  assign n537 = x24 & x82 ;
  assign n538 = n487 & n537 ;
  assign n539 = n491 & n538 ;
  assign n540 = n536 & n539 ;
  assign n541 = ~x129 & ~n540 ;
  assign n544 = ~x45 & ~x49 ;
  assign n545 = ~n257 & n544 ;
  assign n546 = ~n543 & n545 ;
  assign n547 = n254 & n546 ;
  assign n548 = x63 & ~n268 ;
  assign n549 = x82 & n548 ;
  assign n561 = ~x24 & n549 ;
  assign n562 = ~n547 & n561 ;
  assign n560 = ~x24 & ~n548 ;
  assign n563 = n562 ^ n560 ;
  assign n564 = n541 & n563 ;
  assign n565 = ~n559 & n564 ;
  assign n550 = ~n547 & n549 ;
  assign n551 = n550 ^ n548 ;
  assign n552 = n541 & ~n551 ;
  assign n566 = n565 ^ n552 ;
  assign n601 = ~x39 & ~x52 ;
  assign n602 = ~x51 & x116 ;
  assign n603 = n601 & n602 ;
  assign n604 = ~x85 & ~n603 ;
  assign n605 = ~x25 & ~x116 ;
  assign n606 = x26 & ~x27 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = n604 & n607 ;
  assign n592 = ~x85 & ~x96 ;
  assign n593 = x100 & ~x110 ;
  assign n594 = n592 & n593 ;
  assign n590 = x85 & x100 ;
  assign n591 = x116 & n590 ;
  assign n595 = n594 ^ n591 ;
  assign n596 = x85 & ~x116 ;
  assign n597 = x25 & n596 ;
  assign n598 = ~n595 & ~n597 ;
  assign n599 = ~x26 & ~x27 ;
  assign n600 = ~n598 & n599 ;
  assign n609 = n608 ^ n600 ;
  assign n576 = ~x51 & ~x52 ;
  assign n577 = ~x39 & n576 ;
  assign n578 = x27 & ~n577 ;
  assign n579 = x95 & x100 ;
  assign n580 = n579 ^ x95 ;
  assign n581 = n580 ^ x100 ;
  assign n582 = ~x97 & ~x110 ;
  assign n583 = ~n581 & n582 ;
  assign n584 = n583 ^ x110 ;
  assign n585 = x25 & n584 ;
  assign n586 = ~n578 & n585 ;
  assign n587 = ~x26 & ~x85 ;
  assign n613 = n586 & n587 ;
  assign n614 = ~n609 & n613 ;
  assign n615 = n614 ^ n609 ;
  assign n588 = x27 & n587 ;
  assign n589 = ~n586 & n588 ;
  assign n569 = x25 & ~x116 ;
  assign n610 = ~n569 & ~n603 ;
  assign n611 = ~n609 & ~n610 ;
  assign n612 = n589 & n611 ;
  assign n616 = n615 ^ n612 ;
  assign n567 = ~x53 & ~x58 ;
  assign n568 = ~x27 & ~x85 ;
  assign n570 = ~x26 & n569 ;
  assign n571 = n568 & n570 ;
  assign n572 = ~n567 & ~n571 ;
  assign n573 = n204 & ~n572 ;
  assign n574 = x58 ^ x53 ;
  assign n617 = ~x53 & ~n574 ;
  assign n618 = n573 & n617 ;
  assign n619 = n616 & n618 ;
  assign n575 = n573 & n574 ;
  assign n620 = n619 ^ n575 ;
  assign n621 = x26 & ~x85 ;
  assign n622 = ~n603 & n621 ;
  assign n623 = x26 & x116 ;
  assign n624 = n595 & ~n623 ;
  assign n625 = ~n622 & ~n624 ;
  assign n626 = ~x27 & ~x53 ;
  assign n627 = ~x58 & n626 ;
  assign n628 = n204 & n627 ;
  assign n629 = ~n625 & n628 ;
  assign n630 = x27 & n604 ;
  assign n631 = x85 & x116 ;
  assign n632 = ~x85 & ~x110 ;
  assign n633 = x95 & ~x96 ;
  assign n634 = n632 & n633 ;
  assign n635 = ~n631 & ~n634 ;
  assign n636 = ~x27 & ~x100 ;
  assign n637 = ~n635 & n636 ;
  assign n638 = ~n630 & ~n637 ;
  assign n639 = ~x26 & n204 ;
  assign n640 = n567 & n639 ;
  assign n641 = ~n638 & n640 ;
  assign n682 = x26 & x53 ;
  assign n683 = n682 ^ x26 ;
  assign n684 = n683 ^ x53 ;
  assign n685 = x85 & ~n684 ;
  assign n686 = n685 ^ n684 ;
  assign n687 = ~x27 & x28 ;
  assign n688 = ~x116 & n687 ;
  assign n689 = x58 & n688 ;
  assign n690 = ~n686 & n689 ;
  assign n697 = x58 & n204 ;
  assign n698 = ~n690 & n697 ;
  assign n699 = n698 ^ n204 ;
  assign n642 = ~x51 & n601 ;
  assign n643 = n623 & n642 ;
  assign n649 = n568 & n643 ;
  assign n650 = n649 ^ x85 ;
  assign n644 = ~x26 & ~x100 ;
  assign n645 = ~x110 & n644 ;
  assign n646 = n568 & n633 ;
  assign n647 = n645 & n646 ;
  assign n648 = ~n643 & n647 ;
  assign n651 = n650 ^ n648 ;
  assign n652 = ~x26 & x116 ;
  assign n653 = n578 & n652 ;
  assign n654 = ~n651 & n653 ;
  assign n655 = n654 ^ n651 ;
  assign n658 = ~x27 & ~x39 ;
  assign n659 = n576 & n658 ;
  assign n660 = n659 ^ x26 ;
  assign n656 = ~x26 & ~x39 ;
  assign n657 = n576 & n656 ;
  assign n661 = n660 ^ n657 ;
  assign n662 = n584 & ~n661 ;
  assign n663 = x27 ^ x26 ;
  assign n664 = ~x116 & n663 ;
  assign n665 = x28 & ~n664 ;
  assign n666 = ~n662 & n665 ;
  assign n667 = n666 ^ x28 ;
  assign n668 = x100 & x116 ;
  assign n669 = ~x28 & ~x116 ;
  assign n670 = n599 & ~n669 ;
  assign n671 = ~n668 & n670 ;
  assign n677 = ~x53 & n671 ;
  assign n678 = ~n667 & n677 ;
  assign n679 = ~n655 & n678 ;
  assign n680 = n679 ^ n677 ;
  assign n672 = ~x53 & ~x85 ;
  assign n673 = ~n671 & n672 ;
  assign n674 = ~n667 & n673 ;
  assign n675 = ~n655 & n674 ;
  assign n676 = n675 ^ n673 ;
  assign n681 = n680 ^ n676 ;
  assign n691 = ~x58 & n204 ;
  assign n692 = x53 & n587 ;
  assign n693 = n688 & n692 ;
  assign n694 = n691 & ~n693 ;
  assign n695 = ~n690 & n694 ;
  assign n696 = ~n681 & n695 ;
  assign n700 = n699 ^ n696 ;
  assign n701 = x29 & ~x116 ;
  assign n724 = x85 & n701 ;
  assign n725 = n627 & n724 ;
  assign n731 = ~x26 & x85 ;
  assign n732 = ~n725 & n731 ;
  assign n733 = n732 ^ x26 ;
  assign n710 = x29 & x110 ;
  assign n705 = ~x96 & ~x110 ;
  assign n706 = x97 & ~n705 ;
  assign n707 = x29 & ~x110 ;
  assign n708 = ~n581 & n707 ;
  assign n709 = ~n706 & n708 ;
  assign n711 = n710 ^ n709 ;
  assign n712 = ~x58 & x97 ;
  assign n713 = ~n581 & n712 ;
  assign n714 = ~n706 & n713 ;
  assign n715 = n714 ^ x58 ;
  assign n716 = ~n711 & ~n715 ;
  assign n717 = x97 & x116 ;
  assign n718 = x58 & ~n701 ;
  assign n719 = ~n717 & n718 ;
  assign n702 = x53 & ~x58 ;
  assign n703 = n701 & n702 ;
  assign n720 = n626 & ~n703 ;
  assign n721 = ~n719 & n720 ;
  assign n722 = ~n716 & n721 ;
  assign n704 = ~x27 & n703 ;
  assign n723 = n722 ^ n704 ;
  assign n726 = x27 & n567 ;
  assign n727 = n701 & n726 ;
  assign n728 = n587 & ~n727 ;
  assign n729 = ~n725 & n728 ;
  assign n730 = ~n723 & n729 ;
  assign n734 = n733 ^ n730 ;
  assign n735 = ~x85 & n567 ;
  assign n736 = n606 & n735 ;
  assign n737 = n701 & n736 ;
  assign n738 = n204 & ~n737 ;
  assign n739 = n734 & n738 ;
  assign n740 = n739 ^ n204 ;
  assign n741 = ~x30 & ~x109 ;
  assign n742 = ~x60 & x109 ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = ~x106 & ~n743 ;
  assign n745 = ~x88 & x106 ;
  assign n746 = ~x129 & ~n745 ;
  assign n747 = ~n744 & n746 ;
  assign n748 = ~x31 & ~x109 ;
  assign n749 = ~x30 & x109 ;
  assign n750 = ~n748 & ~n749 ;
  assign n751 = ~x106 & ~n750 ;
  assign n752 = ~x89 & x106 ;
  assign n753 = ~x129 & ~n752 ;
  assign n754 = ~n751 & n753 ;
  assign n755 = ~x32 & ~x109 ;
  assign n756 = ~x31 & x109 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = ~x106 & ~n757 ;
  assign n759 = ~x99 & x106 ;
  assign n760 = ~x129 & ~n759 ;
  assign n761 = ~n758 & n760 ;
  assign n762 = ~x33 & ~x109 ;
  assign n763 = ~x32 & x109 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = ~x106 & ~n764 ;
  assign n766 = ~x90 & x106 ;
  assign n767 = ~x129 & ~n766 ;
  assign n768 = ~n765 & n767 ;
  assign n769 = ~x34 & ~x109 ;
  assign n770 = ~x33 & x109 ;
  assign n771 = ~n769 & ~n770 ;
  assign n772 = ~x106 & ~n771 ;
  assign n773 = ~x91 & x106 ;
  assign n774 = ~x129 & ~n773 ;
  assign n775 = ~n772 & n774 ;
  assign n776 = ~x35 & ~x109 ;
  assign n777 = ~x34 & x109 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = ~x106 & ~n778 ;
  assign n780 = ~x92 & x106 ;
  assign n781 = ~x129 & ~n780 ;
  assign n782 = ~n779 & n781 ;
  assign n783 = ~x36 & ~x109 ;
  assign n784 = ~x35 & x109 ;
  assign n785 = ~n783 & ~n784 ;
  assign n786 = ~x106 & ~n785 ;
  assign n787 = ~x98 & x106 ;
  assign n788 = ~x129 & ~n787 ;
  assign n789 = ~n786 & n788 ;
  assign n790 = ~x37 & ~x109 ;
  assign n791 = ~x36 & x109 ;
  assign n792 = ~n790 & ~n791 ;
  assign n793 = ~x106 & ~n792 ;
  assign n794 = ~x93 & x106 ;
  assign n795 = ~x129 & ~n794 ;
  assign n796 = ~n793 & n795 ;
  assign n804 = x82 & ~n282 ;
  assign n808 = ~x38 & n804 ;
  assign n797 = ~x45 & ~x50 ;
  assign n798 = ~n265 & n797 ;
  assign n799 = ~n543 & n798 ;
  assign n800 = x82 & n275 ;
  assign n801 = n418 & n800 ;
  assign n802 = n799 & n801 ;
  assign n803 = n802 ^ x82 ;
  assign n805 = ~x38 & n268 ;
  assign n806 = ~n804 & n805 ;
  assign n807 = ~n803 & n806 ;
  assign n809 = n808 ^ n807 ;
  assign n817 = ~x45 & ~x48 ;
  assign n818 = ~n265 & n817 ;
  assign n819 = ~n543 & n818 ;
  assign n820 = n275 & n277 ;
  assign n821 = ~x40 & ~x50 ;
  assign n822 = ~n252 & n821 ;
  assign n823 = n820 & n822 ;
  assign n824 = n819 & n823 ;
  assign n810 = ~x44 & x82 ;
  assign n811 = ~x40 & ~x42 ;
  assign n812 = x38 & n811 ;
  assign n813 = n810 & n812 ;
  assign n814 = x74 & ~n268 ;
  assign n825 = n445 & n814 ;
  assign n826 = ~n813 & n825 ;
  assign n827 = ~n824 & n826 ;
  assign n815 = ~x129 & ~n814 ;
  assign n816 = ~n813 & n815 ;
  assign n828 = n827 ^ n816 ;
  assign n829 = ~n809 & n828 ;
  assign n830 = x109 & n576 ;
  assign n831 = x39 & ~n830 ;
  assign n832 = ~x51 & x109 ;
  assign n833 = n601 & n832 ;
  assign n834 = ~x106 & ~n833 ;
  assign n835 = ~n831 & n834 ;
  assign n836 = ~x129 & ~n835 ;
  assign n839 = x82 & n252 ;
  assign n843 = ~x40 & n839 ;
  assign n837 = n267 & n280 ;
  assign n838 = n837 ^ x82 ;
  assign n840 = ~x40 & n268 ;
  assign n841 = ~n839 & n840 ;
  assign n842 = ~n838 & n841 ;
  assign n844 = n843 ^ n842 ;
  assign n845 = ~x42 & n810 ;
  assign n846 = x40 & n845 ;
  assign n847 = ~x129 & ~n846 ;
  assign n848 = ~n844 & n847 ;
  assign n860 = x73 & ~n268 ;
  assign n864 = n848 & ~n860 ;
  assign n849 = x46 & ~n244 ;
  assign n850 = n849 ^ n244 ;
  assign n851 = ~n249 & ~n850 ;
  assign n852 = ~n257 & ~n261 ;
  assign n853 = x2 & x45 ;
  assign n854 = n853 ^ x2 ;
  assign n855 = n854 ^ x45 ;
  assign n856 = ~n265 & ~n855 ;
  assign n857 = n852 & n856 ;
  assign n858 = n851 & n857 ;
  assign n859 = ~n252 & n858 ;
  assign n861 = x82 & n860 ;
  assign n862 = ~n859 & n861 ;
  assign n863 = n848 & n862 ;
  assign n865 = n864 ^ n863 ;
  assign n866 = x82 & n268 ;
  assign n867 = n279 & n866 ;
  assign n868 = n274 & n867 ;
  assign n869 = n868 ^ n439 ;
  assign n873 = ~x41 & n869 ;
  assign n870 = ~x41 & x82 ;
  assign n871 = ~n556 & n870 ;
  assign n872 = ~n869 & n871 ;
  assign n874 = n873 ^ n872 ;
  assign n875 = x41 & n845 ;
  assign n876 = n246 & n875 ;
  assign n877 = ~x129 & ~n876 ;
  assign n878 = ~n874 & n877 ;
  assign n881 = x76 & ~n268 ;
  assign n885 = n878 & ~n881 ;
  assign n879 = n274 & n279 ;
  assign n880 = n492 & n879 ;
  assign n882 = x82 & n881 ;
  assign n883 = ~n880 & n882 ;
  assign n884 = n878 & n883 ;
  assign n886 = n885 ^ n884 ;
  assign n902 = ~n249 & n811 ;
  assign n903 = ~n850 & n902 ;
  assign n904 = n857 & n903 ;
  assign n892 = x44 & x82 ;
  assign n896 = ~x42 & n892 ;
  assign n887 = ~x40 & x82 ;
  assign n888 = ~n249 & n887 ;
  assign n889 = ~n850 & n888 ;
  assign n890 = n857 & n889 ;
  assign n891 = n890 ^ x82 ;
  assign n893 = ~x42 & n268 ;
  assign n894 = ~n892 & n893 ;
  assign n895 = ~n891 & n894 ;
  assign n897 = n896 ^ n895 ;
  assign n898 = x42 & n810 ;
  assign n899 = ~x129 & ~n898 ;
  assign n905 = x72 & ~n269 ;
  assign n906 = n899 & n905 ;
  assign n907 = ~n897 & n906 ;
  assign n908 = ~n904 & n907 ;
  assign n900 = ~x72 & n899 ;
  assign n901 = ~n897 & n900 ;
  assign n909 = n908 ^ n901 ;
  assign n910 = ~n423 & n426 ;
  assign n911 = x82 & ~n425 ;
  assign n912 = n910 & n911 ;
  assign n913 = n912 ^ x82 ;
  assign n914 = n268 & n913 ;
  assign n915 = n914 ^ n268 ;
  assign n916 = x82 & ~n415 ;
  assign n917 = ~x43 & ~n916 ;
  assign n918 = ~n915 & n917 ;
  assign n919 = n918 ^ x43 ;
  assign n924 = ~n252 & n887 ;
  assign n925 = n276 & n924 ;
  assign n926 = n857 & n925 ;
  assign n927 = n926 ^ x82 ;
  assign n920 = n810 & n811 ;
  assign n921 = n276 & n920 ;
  assign n928 = x77 & ~n268 ;
  assign n934 = ~x129 & n928 ;
  assign n935 = ~n921 & n934 ;
  assign n936 = ~n927 & n935 ;
  assign n933 = ~x129 & ~n921 ;
  assign n937 = n936 ^ n933 ;
  assign n922 = ~x43 & ~x129 ;
  assign n929 = n922 & n928 ;
  assign n930 = n921 & n929 ;
  assign n931 = ~n927 & n930 ;
  assign n923 = n921 & n922 ;
  assign n932 = n931 ^ n923 ;
  assign n938 = n937 ^ n932 ;
  assign n939 = ~n919 & n938 ;
  assign n940 = n939 ^ n938 ;
  assign n941 = ~x67 & ~n268 ;
  assign n942 = x44 & n268 ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = ~x129 & ~n892 ;
  assign n948 = ~n943 & n944 ;
  assign n945 = x82 & n944 ;
  assign n946 = n943 & n945 ;
  assign n947 = ~n904 & n946 ;
  assign n949 = n948 ^ n947 ;
  assign n950 = x50 & n491 ;
  assign n951 = n950 ^ n491 ;
  assign n952 = n801 & n951 ;
  assign n953 = n952 ^ x82 ;
  assign n954 = n268 & n426 ;
  assign n955 = ~n265 & n496 ;
  assign n956 = n954 & n955 ;
  assign n957 = n956 ^ n439 ;
  assign n958 = ~x45 & ~n957 ;
  assign n959 = ~n953 & n958 ;
  assign n960 = n959 ^ x45 ;
  assign n961 = ~n257 & n426 ;
  assign n962 = ~n423 & n961 ;
  assign n963 = n254 & n962 ;
  assign n964 = x68 & ~n268 ;
  assign n965 = x82 & n964 ;
  assign n966 = ~n963 & n965 ;
  assign n967 = n966 ^ n964 ;
  assign n968 = n275 & n418 ;
  assign n969 = x45 & x82 ;
  assign n970 = ~x50 & ~x129 ;
  assign n971 = n969 & n970 ;
  assign n972 = n491 & n971 ;
  assign n973 = n968 & n972 ;
  assign n974 = n973 ^ x129 ;
  assign n975 = ~n967 & ~n974 ;
  assign n976 = n960 & n975 ;
  assign n977 = ~x75 & n269 ;
  assign n978 = x82 & n951 ;
  assign n979 = x46 & ~n269 ;
  assign n980 = ~n978 & n979 ;
  assign n981 = ~n977 & ~n980 ;
  assign n982 = x82 & ~n249 ;
  assign n983 = n857 & n982 ;
  assign n984 = n983 ^ x82 ;
  assign n985 = ~x75 & ~n268 ;
  assign n986 = n492 & ~n985 ;
  assign n987 = ~n984 & n986 ;
  assign n988 = n987 ^ n492 ;
  assign n989 = ~x129 & ~n988 ;
  assign n990 = n981 & n989 ;
  assign n991 = n990 ^ x129 ;
  assign n993 = n268 & n819 ;
  assign n992 = n439 & ~n819 ;
  assign n994 = n993 ^ n992 ;
  assign n998 = ~x47 & n994 ;
  assign n995 = ~x47 & x82 ;
  assign n996 = ~n254 & n995 ;
  assign n997 = ~n994 & n996 ;
  assign n999 = n998 ^ n997 ;
  assign n1000 = ~x43 & x47 ;
  assign n1001 = n921 & n1000 ;
  assign n1002 = ~x129 & ~n1001 ;
  assign n1003 = ~n999 & n1002 ;
  assign n1005 = x64 & ~n268 ;
  assign n1009 = n1003 & ~n1005 ;
  assign n1004 = n254 & n819 ;
  assign n1006 = x82 & n1005 ;
  assign n1007 = ~n1004 & n1006 ;
  assign n1008 = n1003 & n1007 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1013 = ~x47 & n254 ;
  assign n1014 = ~n417 & ~n543 ;
  assign n1011 = x62 & ~n268 ;
  assign n1015 = x82 & n1011 ;
  assign n1016 = n1014 & n1015 ;
  assign n1017 = n1013 & n1016 ;
  assign n1012 = ~x82 & n1011 ;
  assign n1018 = n1017 ^ n1012 ;
  assign n1019 = x82 & n820 ;
  assign n1020 = n951 & n1019 ;
  assign n1021 = n1020 ^ x82 ;
  assign n1022 = ~x24 & ~x45 ;
  assign n1023 = ~x49 & x82 ;
  assign n1024 = n1022 & n1023 ;
  assign n1025 = ~n543 & n1024 ;
  assign n1026 = n1025 ^ x82 ;
  assign n1033 = x48 & n268 ;
  assign n1034 = ~n1026 & n1033 ;
  assign n1035 = ~n1021 & n1034 ;
  assign n1032 = x48 & ~n1021 ;
  assign n1036 = n1035 ^ n1032 ;
  assign n1037 = n1036 ^ x48 ;
  assign n1027 = n268 & n1026 ;
  assign n1028 = n1027 ^ n268 ;
  assign n1029 = n1021 & n1028 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1031 = n1030 ^ n1021 ;
  assign n1038 = n1037 ^ n1031 ;
  assign n1039 = x48 & n277 ;
  assign n1040 = n921 & n1039 ;
  assign n1041 = ~x129 & ~n1040 ;
  assign n1042 = n1038 & n1041 ;
  assign n1043 = n1042 ^ n1041 ;
  assign n1044 = n1018 & n1043 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n1065 = ~x69 & ~n268 ;
  assign n1061 = n487 & ~n490 ;
  assign n1062 = n435 & n1061 ;
  assign n1063 = n494 & n1062 ;
  assign n1064 = n1063 ^ x82 ;
  assign n1066 = n1065 ^ n1064 ;
  assign n1067 = x49 & n439 ;
  assign n1068 = n1067 ^ n1065 ;
  assign n1069 = n1067 & n1068 ;
  assign n1070 = n1069 ^ n1067 ;
  assign n1071 = n1070 ^ n1064 ;
  assign n1072 = ~n1066 & ~n1071 ;
  assign n1073 = n1072 ^ n1069 ;
  assign n1074 = n1073 ^ n1064 ;
  assign n1046 = n495 & ~n543 ;
  assign n1047 = n1046 ^ n495 ;
  assign n1048 = x24 & x40 ;
  assign n1049 = n1048 ^ x24 ;
  assign n1050 = n1049 ^ x40 ;
  assign n1051 = ~n252 & ~n1050 ;
  assign n1052 = ~n850 & n1051 ;
  assign n1053 = ~n249 & ~n257 ;
  assign n1054 = ~x45 & x49 ;
  assign n1055 = n1053 & n1054 ;
  assign n1056 = n1052 & n1055 ;
  assign n1057 = n1056 ^ x49 ;
  assign n1058 = x82 & ~n1057 ;
  assign n1059 = ~n1047 & n1058 ;
  assign n1060 = n1059 ^ x82 ;
  assign n1075 = n1074 ^ n1060 ;
  assign n1076 = n1074 ^ x129 ;
  assign n1077 = x129 & n1076 ;
  assign n1078 = n1077 ^ x129 ;
  assign n1079 = n1078 ^ n1060 ;
  assign n1080 = ~n1075 & ~n1079 ;
  assign n1081 = n1080 ^ n1077 ;
  assign n1082 = n1081 ^ n1060 ;
  assign n1096 = ~x50 & n820 ;
  assign n1097 = n819 & n1096 ;
  assign n1098 = x82 & ~n1097 ;
  assign n1086 = x82 & ~n491 ;
  assign n1090 = ~x50 & n1086 ;
  assign n1083 = n279 & n800 ;
  assign n1084 = n274 & n1083 ;
  assign n1085 = n1084 ^ x82 ;
  assign n1087 = ~x50 & n268 ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = ~n1085 & n1088 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1092 = x50 & x82 ;
  assign n1093 = n491 & n1092 ;
  assign n1094 = ~x129 & ~n1093 ;
  assign n1099 = x66 & ~n268 ;
  assign n1100 = n1094 & n1099 ;
  assign n1101 = ~n1091 & n1100 ;
  assign n1102 = ~n1098 & n1101 ;
  assign n1095 = ~n1091 & n1094 ;
  assign n1103 = n1102 ^ n1095 ;
  assign n1104 = x51 & ~x109 ;
  assign n1105 = ~x106 & ~n832 ;
  assign n1106 = ~n1104 & n1105 ;
  assign n1107 = ~x129 & ~n1106 ;
  assign n1108 = x52 & ~n832 ;
  assign n1109 = ~x106 & ~n830 ;
  assign n1110 = ~n1108 & n1109 ;
  assign n1111 = ~x129 & ~n1110 ;
  assign n1112 = ~x116 & n702 ;
  assign n1113 = ~x53 & x97 ;
  assign n1114 = x58 & x116 ;
  assign n1115 = ~x58 & ~n581 ;
  assign n1116 = n705 & n1115 ;
  assign n1117 = ~n1114 & ~n1116 ;
  assign n1118 = n1113 & ~n1117 ;
  assign n1119 = ~n1112 & ~n1118 ;
  assign n1120 = n568 & n639 ;
  assign n1121 = ~n1119 & n1120 ;
  assign n1122 = ~n268 & n910 ;
  assign n1123 = n557 & n1122 ;
  assign n1124 = ~x129 & ~n269 ;
  assign n1125 = ~n1123 & n1124 ;
  assign n1126 = ~x123 & ~x129 ;
  assign n1127 = x114 & ~x122 ;
  assign n1128 = n1126 & n1127 ;
  assign n1138 = x37 & ~x58 ;
  assign n1139 = ~x116 & n1138 ;
  assign n1135 = x26 & ~x58 ;
  assign n1136 = x94 & x116 ;
  assign n1137 = n1135 & n1136 ;
  assign n1140 = n1139 ^ n1137 ;
  assign n1131 = ~x26 & x58 ;
  assign n1132 = ~x94 & ~x116 ;
  assign n1133 = n1131 & n1132 ;
  assign n1134 = n1133 ^ n1131 ;
  assign n1141 = n1140 ^ n1134 ;
  assign n1129 = ~x26 & x37 ;
  assign n1144 = n567 & n1129 ;
  assign n1145 = n1141 & n1144 ;
  assign n1143 = ~x58 & n1129 ;
  assign n1146 = n1145 ^ n1143 ;
  assign n1142 = ~x53 & n1141 ;
  assign n1147 = n1146 ^ n1142 ;
  assign n1154 = n568 & n1147 ;
  assign n1152 = x85 & n567 ;
  assign n1153 = n1129 & n1152 ;
  assign n1155 = n1154 ^ n1153 ;
  assign n1148 = n568 & n1129 ;
  assign n1149 = n567 & n1148 ;
  assign n1150 = ~n1147 & n1149 ;
  assign n1130 = n726 & n1129 ;
  assign n1151 = n1150 ^ n1130 ;
  assign n1156 = n1155 ^ n1151 ;
  assign n1157 = n204 & n1156 ;
  assign n1175 = x60 & n1114 ;
  assign n1176 = ~n686 & n1175 ;
  assign n1158 = ~x85 & ~x116 ;
  assign n1159 = ~n684 & n1158 ;
  assign n1162 = x85 ^ x53 ;
  assign n1163 = n1162 ^ x85 ;
  assign n1160 = x85 ^ x26 ;
  assign n1161 = n1160 ^ x85 ;
  assign n1164 = n1163 ^ n1161 ;
  assign n1165 = n1163 ^ x85 ;
  assign n1166 = n1164 & n1165 ;
  assign n1167 = n1166 ^ n1163 ;
  assign n1168 = ~x58 & n1167 ;
  assign n1169 = n1168 ^ x58 ;
  assign n1170 = n1159 & ~n1169 ;
  assign n1171 = n1170 ^ n1159 ;
  assign n1172 = n1171 ^ n1169 ;
  assign n1173 = x57 & n1172 ;
  assign n1174 = n1173 ^ x57 ;
  assign n1177 = n1176 ^ n1174 ;
  assign n1178 = n1176 ^ x27 ;
  assign n1179 = x27 & ~n1178 ;
  assign n1180 = n1179 ^ x27 ;
  assign n1181 = n1180 ^ n1174 ;
  assign n1182 = n1177 & ~n1181 ;
  assign n1183 = n1182 ^ n1179 ;
  assign n1184 = n1183 ^ n1174 ;
  assign n1185 = x57 & ~x58 ;
  assign n1186 = ~n686 & n1185 ;
  assign n1187 = n1184 & n1186 ;
  assign n1188 = n1187 ^ n1184 ;
  assign n1189 = n1188 ^ n1186 ;
  assign n1190 = n204 & ~n1189 ;
  assign n1191 = n1190 ^ n204 ;
  assign n1192 = x58 & ~x116 ;
  assign n1193 = n599 & n1192 ;
  assign n1194 = ~x58 & n663 ;
  assign n1195 = n603 & n1194 ;
  assign n1196 = ~n1193 & ~n1195 ;
  assign n1197 = n204 & n672 ;
  assign n1198 = ~n1196 & n1197 ;
  assign n1199 = x59 & ~x116 ;
  assign n1215 = n735 & n1199 ;
  assign n1216 = n204 & n663 ;
  assign n1217 = n1215 & n1216 ;
  assign n1218 = n1217 ^ n204 ;
  assign n1203 = x96 ^ x59 ;
  assign n1204 = n567 & n1203 ;
  assign n1205 = n584 & n1204 ;
  assign n1202 = x96 & n567 ;
  assign n1206 = n1205 ^ n1202 ;
  assign n1201 = n574 & n1199 ;
  assign n1207 = n1206 ^ n1201 ;
  assign n1208 = n1207 ^ x85 ;
  assign n1209 = n1207 & ~n1208 ;
  assign n1200 = n1152 & n1199 ;
  assign n1210 = n1209 ^ n1200 ;
  assign n1211 = n1210 ^ n1207 ;
  assign n1212 = ~x27 & ~n663 ;
  assign n1213 = n204 & n1212 ;
  assign n1214 = n1211 & n1213 ;
  assign n1219 = n1218 ^ n1214 ;
  assign n1220 = n1219 ^ n204 ;
  assign n1221 = ~x117 & ~x122 ;
  assign n1222 = x60 & ~n1221 ;
  assign n1223 = x123 & n1221 ;
  assign n1224 = ~n1222 & ~n1223 ;
  assign n1225 = ~x114 & ~x122 ;
  assign n1226 = x123 & ~x129 ;
  assign n1227 = n1225 & n1226 ;
  assign n1228 = x136 & ~x137 ;
  assign n1229 = x131 & x132 ;
  assign n1230 = x133 & n1229 ;
  assign n1231 = ~x138 & n1230 ;
  assign n1232 = n1228 & n1231 ;
  assign n1233 = x140 & n1232 ;
  assign n1234 = ~x62 & ~n1232 ;
  assign n1235 = ~x129 & ~n1234 ;
  assign n1236 = ~n1233 & n1235 ;
  assign n1237 = x142 & n1232 ;
  assign n1238 = ~x63 & ~n1232 ;
  assign n1239 = ~x129 & ~n1238 ;
  assign n1240 = ~n1237 & n1239 ;
  assign n1241 = x139 & n1232 ;
  assign n1242 = ~x64 & ~n1232 ;
  assign n1243 = ~x129 & ~n1242 ;
  assign n1244 = ~n1241 & n1243 ;
  assign n1245 = x146 & n1232 ;
  assign n1246 = ~x65 & ~n1232 ;
  assign n1247 = ~x129 & ~n1246 ;
  assign n1248 = ~n1245 & n1247 ;
  assign n1249 = ~x136 & ~x137 ;
  assign n1250 = n1231 & n1249 ;
  assign n1251 = x143 & n1250 ;
  assign n1252 = ~x66 & ~n1250 ;
  assign n1253 = ~x129 & ~n1252 ;
  assign n1254 = ~n1251 & n1253 ;
  assign n1255 = x139 & n1250 ;
  assign n1256 = ~x67 & ~n1250 ;
  assign n1257 = ~x129 & ~n1256 ;
  assign n1258 = ~n1255 & n1257 ;
  assign n1259 = x141 & n1232 ;
  assign n1260 = ~x68 & ~n1232 ;
  assign n1261 = ~x129 & ~n1260 ;
  assign n1262 = ~n1259 & n1261 ;
  assign n1263 = x143 & n1232 ;
  assign n1264 = ~x69 & ~n1232 ;
  assign n1265 = ~x129 & ~n1264 ;
  assign n1266 = ~n1263 & n1265 ;
  assign n1267 = x144 & n1232 ;
  assign n1268 = ~x70 & ~n1232 ;
  assign n1269 = ~x129 & ~n1268 ;
  assign n1270 = ~n1267 & n1269 ;
  assign n1271 = x145 & n1232 ;
  assign n1272 = ~x71 & ~n1232 ;
  assign n1273 = ~x129 & ~n1272 ;
  assign n1274 = ~n1271 & n1273 ;
  assign n1275 = x140 & n1250 ;
  assign n1276 = ~x72 & ~n1250 ;
  assign n1277 = ~x129 & ~n1276 ;
  assign n1278 = ~n1275 & n1277 ;
  assign n1279 = x141 & n1250 ;
  assign n1280 = ~x73 & ~n1250 ;
  assign n1281 = ~x129 & ~n1280 ;
  assign n1282 = ~n1279 & n1281 ;
  assign n1283 = x142 & n1250 ;
  assign n1284 = ~x74 & ~n1250 ;
  assign n1285 = ~x129 & ~n1284 ;
  assign n1286 = ~n1283 & n1285 ;
  assign n1287 = x144 & n1250 ;
  assign n1288 = ~x75 & ~n1250 ;
  assign n1289 = ~x129 & ~n1288 ;
  assign n1290 = ~n1287 & n1289 ;
  assign n1291 = x145 & n1250 ;
  assign n1292 = ~x76 & ~n1250 ;
  assign n1293 = ~x129 & ~n1292 ;
  assign n1294 = ~n1291 & n1293 ;
  assign n1295 = x146 & n1250 ;
  assign n1296 = ~x77 & ~n1250 ;
  assign n1297 = ~x129 & ~n1296 ;
  assign n1298 = ~n1295 & n1297 ;
  assign n1299 = ~x136 & x137 ;
  assign n1300 = n1231 & n1299 ;
  assign n1301 = ~x142 & n1300 ;
  assign n1302 = ~x78 & ~n1300 ;
  assign n1303 = ~x129 & ~n1302 ;
  assign n1304 = ~n1301 & n1303 ;
  assign n1305 = ~x143 & n1300 ;
  assign n1306 = ~x79 & ~n1300 ;
  assign n1307 = ~x129 & ~n1306 ;
  assign n1308 = ~n1305 & n1307 ;
  assign n1309 = ~x144 & n1300 ;
  assign n1310 = ~x80 & ~n1300 ;
  assign n1311 = ~x129 & ~n1310 ;
  assign n1312 = ~n1309 & n1311 ;
  assign n1313 = ~x145 & n1300 ;
  assign n1314 = ~x81 & ~n1300 ;
  assign n1315 = ~x129 & ~n1314 ;
  assign n1316 = ~n1313 & n1315 ;
  assign n1317 = ~x146 & n1300 ;
  assign n1318 = ~x82 & ~n1300 ;
  assign n1319 = ~x129 & ~n1318 ;
  assign n1320 = ~n1317 & n1319 ;
  assign n1321 = x136 & ~x138 ;
  assign n1322 = x31 & n1321 ;
  assign n1323 = x115 & x138 ;
  assign n1324 = ~x87 & ~x138 ;
  assign n1325 = ~x136 & ~n1324 ;
  assign n1326 = ~n1323 & n1325 ;
  assign n1327 = ~n1322 & ~n1326 ;
  assign n1328 = x137 & ~n1327 ;
  assign n1329 = x62 & ~x138 ;
  assign n1330 = ~x89 & x138 ;
  assign n1331 = x136 & ~n1330 ;
  assign n1332 = ~n1329 & n1331 ;
  assign n1333 = x72 & ~x138 ;
  assign n1334 = ~x119 & x138 ;
  assign n1335 = ~x136 & ~n1334 ;
  assign n1336 = ~n1333 & n1335 ;
  assign n1337 = ~n1332 & ~n1336 ;
  assign n1338 = ~x137 & ~n1337 ;
  assign n1339 = ~n1328 & ~n1338 ;
  assign n1340 = ~x141 & n1300 ;
  assign n1341 = ~x84 & ~n1300 ;
  assign n1342 = ~x129 & ~n1341 ;
  assign n1343 = ~n1340 & n1342 ;
  assign n1344 = x97 & ~n581 ;
  assign n1345 = n1344 ^ n581 ;
  assign n1346 = n632 & n1345 ;
  assign n1347 = x96 & n1346 ;
  assign n1348 = ~n596 & ~n1347 ;
  assign n1349 = n627 & n639 ;
  assign n1350 = ~n1348 & n1349 ;
  assign n1351 = ~x139 & n1300 ;
  assign n1352 = ~x86 & ~n1300 ;
  assign n1353 = ~x129 & ~n1352 ;
  assign n1354 = ~n1351 & n1353 ;
  assign n1355 = ~x140 & n1300 ;
  assign n1356 = ~x87 & ~n1300 ;
  assign n1357 = ~x129 & ~n1356 ;
  assign n1358 = ~n1355 & n1357 ;
  assign n1359 = x137 & n1321 ;
  assign n1360 = n1230 & n1359 ;
  assign n1361 = ~x139 & n1360 ;
  assign n1362 = ~x88 & ~n1360 ;
  assign n1363 = ~x129 & ~n1362 ;
  assign n1364 = ~n1361 & n1363 ;
  assign n1365 = ~x140 & n1360 ;
  assign n1366 = ~x89 & ~n1360 ;
  assign n1367 = ~x129 & ~n1366 ;
  assign n1368 = ~n1365 & n1367 ;
  assign n1369 = ~x142 & n1360 ;
  assign n1370 = ~x90 & ~n1360 ;
  assign n1371 = ~x129 & ~n1370 ;
  assign n1372 = ~n1369 & n1371 ;
  assign n1373 = ~x143 & n1360 ;
  assign n1374 = ~x91 & ~n1360 ;
  assign n1375 = ~x129 & ~n1374 ;
  assign n1376 = ~n1373 & n1375 ;
  assign n1377 = ~x144 & n1360 ;
  assign n1378 = ~x92 & ~n1360 ;
  assign n1379 = ~x129 & ~n1378 ;
  assign n1380 = ~n1377 & n1379 ;
  assign n1381 = ~x146 & n1360 ;
  assign n1382 = ~x93 & ~n1360 ;
  assign n1383 = ~x129 & ~n1382 ;
  assign n1384 = ~n1381 & n1383 ;
  assign n1385 = x82 & x138 ;
  assign n1386 = n1249 & n1385 ;
  assign n1387 = n1230 & n1386 ;
  assign n1388 = ~x142 & n1387 ;
  assign n1389 = ~x94 & ~n1387 ;
  assign n1390 = ~x129 & ~n1389 ;
  assign n1391 = ~n1388 & n1390 ;
  assign n1392 = ~x3 & ~x110 ;
  assign n1393 = ~n1230 & ~n1392 ;
  assign n1394 = ~n1387 & ~n1393 ;
  assign n1395 = x95 & n1394 ;
  assign n1396 = x143 & n1387 ;
  assign n1397 = ~n1395 & ~n1396 ;
  assign n1398 = ~x129 & ~n1397 ;
  assign n1399 = x96 & n1394 ;
  assign n1400 = x146 & n1387 ;
  assign n1401 = ~n1399 & ~n1400 ;
  assign n1402 = ~x129 & ~n1401 ;
  assign n1403 = x97 & n1394 ;
  assign n1404 = x145 & n1387 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~x129 & ~n1405 ;
  assign n1407 = ~x145 & n1360 ;
  assign n1408 = ~x98 & ~n1360 ;
  assign n1409 = ~x129 & ~n1408 ;
  assign n1410 = ~n1407 & n1409 ;
  assign n1411 = ~x141 & n1360 ;
  assign n1412 = ~x99 & ~n1360 ;
  assign n1413 = ~x129 & ~n1412 ;
  assign n1414 = ~n1411 & n1413 ;
  assign n1415 = x100 & n1394 ;
  assign n1416 = x144 & n1387 ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = ~x129 & ~n1417 ;
  assign n1419 = x37 & n1321 ;
  assign n1420 = ~x96 & x138 ;
  assign n1421 = ~x82 & ~x138 ;
  assign n1422 = ~x136 & ~n1421 ;
  assign n1423 = ~n1420 & n1422 ;
  assign n1424 = ~n1419 & ~n1423 ;
  assign n1425 = x137 & ~n1424 ;
  assign n1426 = x65 & ~x138 ;
  assign n1427 = ~x93 & x138 ;
  assign n1428 = x136 & ~n1427 ;
  assign n1429 = ~n1426 & n1428 ;
  assign n1430 = x77 & ~x138 ;
  assign n1431 = ~x124 & x138 ;
  assign n1432 = ~x136 & ~n1431 ;
  assign n1433 = ~n1430 & n1432 ;
  assign n1434 = ~n1429 & ~n1433 ;
  assign n1435 = ~x137 & ~n1434 ;
  assign n1436 = ~n1425 & ~n1435 ;
  assign n1437 = x91 & n1228 ;
  assign n1438 = x95 & n1299 ;
  assign n1439 = ~n1437 & ~n1438 ;
  assign n1440 = x138 & ~n1439 ;
  assign n1441 = ~x34 & x136 ;
  assign n1442 = ~x79 & ~x136 ;
  assign n1443 = x137 & ~n1442 ;
  assign n1444 = ~n1441 & n1443 ;
  assign n1445 = x69 & x136 ;
  assign n1446 = x66 & ~x136 ;
  assign n1447 = ~x137 & ~n1446 ;
  assign n1448 = ~n1445 & n1447 ;
  assign n1449 = ~n1444 & ~n1448 ;
  assign n1450 = ~x138 & ~n1449 ;
  assign n1451 = ~n1440 & ~n1450 ;
  assign n1452 = x90 & n1228 ;
  assign n1453 = x94 & n1299 ;
  assign n1454 = ~n1452 & ~n1453 ;
  assign n1455 = x138 & ~n1454 ;
  assign n1456 = ~x33 & x136 ;
  assign n1457 = ~x78 & ~x136 ;
  assign n1458 = x137 & ~n1457 ;
  assign n1459 = ~n1456 & n1458 ;
  assign n1460 = x63 & x136 ;
  assign n1461 = x74 & ~x136 ;
  assign n1462 = ~x137 & ~n1461 ;
  assign n1463 = ~n1460 & n1462 ;
  assign n1464 = ~n1459 & ~n1463 ;
  assign n1465 = ~x138 & ~n1464 ;
  assign n1466 = ~n1455 & ~n1465 ;
  assign n1467 = x99 & n1228 ;
  assign n1468 = ~x112 & n1299 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = x138 & ~n1469 ;
  assign n1471 = ~x32 & x136 ;
  assign n1472 = ~x84 & ~x136 ;
  assign n1473 = x137 & ~n1472 ;
  assign n1474 = ~n1471 & n1473 ;
  assign n1475 = x68 & x136 ;
  assign n1476 = x73 & ~x136 ;
  assign n1477 = ~x137 & ~n1476 ;
  assign n1478 = ~n1475 & n1477 ;
  assign n1479 = ~n1474 & ~n1478 ;
  assign n1480 = ~x138 & ~n1479 ;
  assign n1481 = ~n1470 & ~n1480 ;
  assign n1482 = x35 & n1321 ;
  assign n1483 = ~x100 & x138 ;
  assign n1484 = ~x80 & ~x138 ;
  assign n1485 = ~x136 & ~n1484 ;
  assign n1486 = ~n1483 & n1485 ;
  assign n1487 = ~n1482 & ~n1486 ;
  assign n1488 = x137 & ~n1487 ;
  assign n1489 = x70 & ~x138 ;
  assign n1490 = ~x92 & x138 ;
  assign n1491 = x136 & ~n1490 ;
  assign n1492 = ~n1489 & n1491 ;
  assign n1493 = x75 & ~x138 ;
  assign n1494 = ~x125 & x138 ;
  assign n1495 = ~x136 & ~n1494 ;
  assign n1496 = ~n1493 & n1495 ;
  assign n1497 = ~n1492 & ~n1496 ;
  assign n1498 = ~x137 & ~n1497 ;
  assign n1499 = ~n1488 & ~n1498 ;
  assign n1500 = ~x26 & n627 ;
  assign n1501 = n1346 & n1500 ;
  assign n1502 = ~n631 & ~n1501 ;
  assign n1503 = n204 & ~n1502 ;
  assign n1504 = x36 & n1321 ;
  assign n1505 = ~x97 & x138 ;
  assign n1506 = ~x81 & ~x138 ;
  assign n1507 = ~x136 & ~n1506 ;
  assign n1508 = ~n1505 & n1507 ;
  assign n1509 = ~n1504 & ~n1508 ;
  assign n1510 = x137 & ~n1509 ;
  assign n1511 = x71 & ~x138 ;
  assign n1512 = ~x98 & x138 ;
  assign n1513 = x136 & ~n1512 ;
  assign n1514 = ~n1511 & n1513 ;
  assign n1515 = x76 & ~x138 ;
  assign n1516 = ~x23 & x138 ;
  assign n1517 = ~x136 & ~n1516 ;
  assign n1518 = ~n1515 & n1517 ;
  assign n1519 = ~n1514 & ~n1518 ;
  assign n1520 = ~x137 & ~n1519 ;
  assign n1521 = ~n1510 & ~n1520 ;
  assign n1522 = x30 & n1321 ;
  assign n1523 = ~x111 & x138 ;
  assign n1524 = ~x86 & ~x138 ;
  assign n1525 = ~x136 & ~n1524 ;
  assign n1526 = ~n1523 & n1525 ;
  assign n1527 = ~n1522 & ~n1526 ;
  assign n1528 = x137 & ~n1527 ;
  assign n1529 = x64 & ~x138 ;
  assign n1530 = ~x88 & x138 ;
  assign n1531 = x136 & ~n1530 ;
  assign n1532 = ~n1529 & n1531 ;
  assign n1533 = x67 & ~x138 ;
  assign n1534 = ~x120 & x138 ;
  assign n1535 = ~x136 & ~n1534 ;
  assign n1536 = ~n1533 & n1535 ;
  assign n1537 = ~n1532 & ~n1536 ;
  assign n1538 = ~x137 & ~n1537 ;
  assign n1539 = ~n1528 & ~n1538 ;
  assign n1540 = ~x26 & n578 ;
  assign n1541 = ~n606 & ~n1540 ;
  assign n1542 = x116 & n204 ;
  assign n1543 = ~n1541 & n1542 ;
  assign n1544 = ~x53 & x58 ;
  assign n1545 = ~x97 & n1544 ;
  assign n1546 = ~n702 & ~n1545 ;
  assign n1547 = n1542 & ~n1546 ;
  assign n1548 = ~x139 & n1386 ;
  assign n1549 = ~x129 & n1230 ;
  assign n1550 = ~x111 & ~n1386 ;
  assign n1551 = n1549 & ~n1550 ;
  assign n1552 = ~n1548 & n1551 ;
  assign n1553 = x112 & ~n1386 ;
  assign n1554 = ~x141 & n1386 ;
  assign n1555 = n1549 & ~n1554 ;
  assign n1556 = ~n1553 & n1555 ;
  assign n1557 = ~x11 & ~x22 ;
  assign n1558 = x54 & n1557 ;
  assign n1559 = ~x54 & x113 ;
  assign n1560 = n204 & ~n1559 ;
  assign n1561 = ~n1558 & n1560 ;
  assign n1562 = x115 & ~n1386 ;
  assign n1563 = ~x140 & n1386 ;
  assign n1564 = n1549 & ~n1563 ;
  assign n1565 = ~n1562 & n1564 ;
  assign n1566 = x54 & n204 ;
  assign n1567 = ~x4 & ~x9 ;
  assign n1568 = n207 & n1567 ;
  assign n1569 = n1566 & ~n1568 ;
  assign n1570 = x122 & ~x129 ;
  assign n1571 = ~x54 & x118 ;
  assign n1572 = x54 & ~x59 ;
  assign n1573 = n397 & n1572 ;
  assign n1574 = ~n1571 & ~n1573 ;
  assign n1575 = ~x129 & ~n1574 ;
  assign n1576 = ~x129 & n581 ;
  assign n1577 = ~x120 & n1392 ;
  assign n1578 = ~x111 & ~x129 ;
  assign n1579 = ~n1577 & n1578 ;
  assign n1580 = x81 & x120 ;
  assign n1581 = ~x129 & n1580 ;
  assign n1582 = ~x129 & ~x134 ;
  assign n1583 = ~x129 & ~x135 ;
  assign n1584 = x57 & ~x129 ;
  assign n1585 = ~x96 & x125 ;
  assign n1586 = ~x3 & ~n1585 ;
  assign n1587 = ~x129 & ~n1586 ;
  assign n1588 = ~x126 & x132 ;
  assign n1589 = x133 & n1588 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n205 ;
  assign y16 = ~n241 ;
  assign y17 = n292 ;
  assign y18 = ~n307 ;
  assign y19 = n323 ;
  assign y20 = n336 ;
  assign y21 = n344 ;
  assign y22 = n351 ;
  assign y23 = n362 ;
  assign y24 = n369 ;
  assign y25 = n379 ;
  assign y26 = n388 ;
  assign y27 = n395 ;
  assign y28 = n406 ;
  assign y29 = n414 ;
  assign y30 = n449 ;
  assign y31 = n457 ;
  assign y32 = n466 ;
  assign y33 = n476 ;
  assign y34 = n485 ;
  assign y35 = n515 ;
  assign y36 = n523 ;
  assign y37 = n532 ;
  assign y38 = n535 ;
  assign y39 = n566 ;
  assign y40 = n620 ;
  assign y41 = n629 ;
  assign y42 = n641 ;
  assign y43 = n700 ;
  assign y44 = n740 ;
  assign y45 = n747 ;
  assign y46 = n754 ;
  assign y47 = n761 ;
  assign y48 = n768 ;
  assign y49 = n775 ;
  assign y50 = n782 ;
  assign y51 = n789 ;
  assign y52 = n796 ;
  assign y53 = n829 ;
  assign y54 = n836 ;
  assign y55 = n865 ;
  assign y56 = n886 ;
  assign y57 = n909 ;
  assign y58 = n940 ;
  assign y59 = n949 ;
  assign y60 = n976 ;
  assign y61 = ~n991 ;
  assign y62 = n1010 ;
  assign y63 = n1045 ;
  assign y64 = n1082 ;
  assign y65 = n1103 ;
  assign y66 = n1107 ;
  assign y67 = n1111 ;
  assign y68 = n1121 ;
  assign y69 = ~n1125 ;
  assign y70 = n1128 ;
  assign y71 = n1157 ;
  assign y72 = n1191 ;
  assign y73 = n1198 ;
  assign y74 = n1220 ;
  assign y75 = ~n1224 ;
  assign y76 = n1227 ;
  assign y77 = ~n1236 ;
  assign y78 = ~n1240 ;
  assign y79 = ~n1244 ;
  assign y80 = ~n1248 ;
  assign y81 = ~n1254 ;
  assign y82 = ~n1258 ;
  assign y83 = ~n1262 ;
  assign y84 = ~n1266 ;
  assign y85 = ~n1270 ;
  assign y86 = ~n1274 ;
  assign y87 = ~n1278 ;
  assign y88 = ~n1282 ;
  assign y89 = ~n1286 ;
  assign y90 = ~n1290 ;
  assign y91 = ~n1294 ;
  assign y92 = ~n1298 ;
  assign y93 = n1304 ;
  assign y94 = n1308 ;
  assign y95 = n1312 ;
  assign y96 = n1316 ;
  assign y97 = n1320 ;
  assign y98 = ~n1339 ;
  assign y99 = n1343 ;
  assign y100 = n1350 ;
  assign y101 = n1354 ;
  assign y102 = n1358 ;
  assign y103 = n1364 ;
  assign y104 = n1368 ;
  assign y105 = n1372 ;
  assign y106 = n1376 ;
  assign y107 = n1380 ;
  assign y108 = n1384 ;
  assign y109 = n1391 ;
  assign y110 = n1398 ;
  assign y111 = n1402 ;
  assign y112 = n1406 ;
  assign y113 = n1410 ;
  assign y114 = n1414 ;
  assign y115 = n1418 ;
  assign y116 = ~n1436 ;
  assign y117 = ~n1451 ;
  assign y118 = ~n1466 ;
  assign y119 = ~n1481 ;
  assign y120 = ~n1499 ;
  assign y121 = n1503 ;
  assign y122 = ~n1521 ;
  assign y123 = ~n1539 ;
  assign y124 = n1543 ;
  assign y125 = n1547 ;
  assign y126 = n1552 ;
  assign y127 = n1556 ;
  assign y128 = n1561 ;
  assign y129 = ~n1126 ;
  assign y130 = n1565 ;
  assign y131 = n1569 ;
  assign y132 = ~n1570 ;
  assign y133 = n1575 ;
  assign y134 = n1576 ;
  assign y135 = n1579 ;
  assign y136 = n1581 ;
  assign y137 = ~n1582 ;
  assign y138 = ~n1583 ;
  assign y139 = n1584 ;
  assign y140 = n1587 ;
  assign y141 = n1589 ;
endmodule
