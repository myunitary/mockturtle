module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 ;
  assign n289 = ~x30 & ~x286 ;
  assign n290 = x30 & x286 ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = ~x29 & ~x285 ;
  assign n293 = x29 & x285 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = n291 & n294 ;
  assign n296 = ~n291 & ~n294 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = ~x31 & ~x287 ;
  assign n299 = x31 & x287 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = ~n297 & ~n300 ;
  assign n302 = n297 & n300 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~x25 & ~x281 ;
  assign n305 = x25 & x281 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = ~n303 & ~n306 ;
  assign n308 = n303 & n306 ;
  assign n309 = ~n307 & ~n308 ;
  assign n310 = ~x27 & ~x283 ;
  assign n311 = x27 & x283 ;
  assign n312 = ~n310 & ~n311 ;
  assign n313 = ~x26 & ~x282 ;
  assign n314 = x26 & x282 ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = ~n312 & ~n315 ;
  assign n317 = n312 & n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~x28 & ~x284 ;
  assign n320 = x28 & x284 ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = ~n318 & ~n321 ;
  assign n323 = n318 & n321 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n309 & ~n324 ;
  assign n326 = ~n307 & ~n325 ;
  assign n327 = ~n295 & ~n302 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = n326 & ~n327 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n317 & ~n323 ;
  assign n332 = n330 & n331 ;
  assign n333 = ~n328 & ~n332 ;
  assign n334 = ~n330 & ~n331 ;
  assign n335 = ~n332 & ~n334 ;
  assign n336 = ~n309 & n324 ;
  assign n337 = ~n325 & ~n336 ;
  assign n338 = ~x17 & ~x273 ;
  assign n339 = x17 & x273 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n337 & ~n340 ;
  assign n342 = ~x23 & ~x279 ;
  assign n343 = x23 & x279 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = ~x22 & ~x278 ;
  assign n346 = x22 & x278 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n344 & ~n347 ;
  assign n349 = n344 & n347 ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = ~x24 & ~x280 ;
  assign n352 = x24 & x280 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = ~n350 & ~n353 ;
  assign n355 = n350 & n353 ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = ~x18 & ~x274 ;
  assign n358 = x18 & x274 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = ~n356 & ~n359 ;
  assign n361 = n356 & n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~x20 & ~x276 ;
  assign n364 = x20 & x276 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = ~x19 & ~x275 ;
  assign n367 = x19 & x275 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = ~n365 & ~n368 ;
  assign n370 = n365 & n368 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = ~x21 & ~x277 ;
  assign n373 = x21 & x277 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = ~n371 & ~n374 ;
  assign n376 = n371 & n374 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = n362 & ~n377 ;
  assign n379 = ~n362 & n377 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n337 & n340 ;
  assign n382 = ~n341 & ~n381 ;
  assign n383 = n380 & n382 ;
  assign n384 = ~n341 & ~n383 ;
  assign n385 = n335 & ~n384 ;
  assign n386 = ~n360 & ~n378 ;
  assign n387 = ~n349 & ~n355 ;
  assign n388 = ~n386 & n387 ;
  assign n389 = n386 & ~n387 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = ~n370 & ~n376 ;
  assign n392 = n390 & n391 ;
  assign n393 = ~n390 & ~n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n335 & n384 ;
  assign n396 = ~n385 & ~n395 ;
  assign n397 = n394 & n396 ;
  assign n398 = ~n385 & ~n397 ;
  assign n399 = ~n333 & ~n398 ;
  assign n400 = n333 & n398 ;
  assign n401 = ~n399 & ~n400 ;
  assign n402 = ~n388 & ~n392 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = ~n399 & ~n403 ;
  assign n405 = ~n401 & n402 ;
  assign n406 = ~n403 & ~n405 ;
  assign n407 = ~n394 & ~n396 ;
  assign n408 = ~n397 & ~n407 ;
  assign n409 = ~n380 & ~n382 ;
  assign n410 = ~n383 & ~n409 ;
  assign n411 = ~x1 & ~x257 ;
  assign n412 = x1 & x257 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = n410 & ~n413 ;
  assign n415 = ~x8 & ~x264 ;
  assign n416 = x8 & x264 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = ~x7 & ~x263 ;
  assign n419 = x7 & x263 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n417 & ~n420 ;
  assign n422 = n417 & n420 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~x9 & ~x265 ;
  assign n425 = x9 & x265 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~n423 & ~n426 ;
  assign n428 = n423 & n426 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = ~x3 & ~x259 ;
  assign n431 = x3 & x259 ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = ~n429 & ~n432 ;
  assign n434 = n429 & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = ~x5 & ~x261 ;
  assign n437 = x5 & x261 ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = ~x4 & ~x260 ;
  assign n440 = x4 & x260 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~n438 & ~n441 ;
  assign n443 = n438 & n441 ;
  assign n444 = ~n442 & ~n443 ;
  assign n445 = ~x6 & ~x262 ;
  assign n446 = x6 & x262 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n444 & ~n447 ;
  assign n449 = n444 & n447 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = n435 & ~n450 ;
  assign n452 = ~n435 & n450 ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = ~x15 & ~x271 ;
  assign n455 = x15 & x271 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = ~x14 & ~x270 ;
  assign n458 = x14 & x270 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = ~n456 & ~n459 ;
  assign n461 = n456 & n459 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~x16 & ~x272 ;
  assign n464 = x16 & x272 ;
  assign n465 = ~n463 & ~n464 ;
  assign n466 = ~n462 & ~n465 ;
  assign n467 = n462 & n465 ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = ~x10 & ~x266 ;
  assign n470 = x10 & x266 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~n468 & ~n471 ;
  assign n473 = n468 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~x12 & ~x268 ;
  assign n476 = x12 & x268 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~x11 & ~x267 ;
  assign n479 = x11 & x267 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = ~n477 & ~n480 ;
  assign n482 = n477 & n480 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = ~x13 & ~x269 ;
  assign n485 = x13 & x269 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~n483 & ~n486 ;
  assign n488 = n483 & n486 ;
  assign n489 = ~n487 & ~n488 ;
  assign n490 = n474 & ~n489 ;
  assign n491 = ~n474 & n489 ;
  assign n492 = ~n490 & ~n491 ;
  assign n493 = ~x2 & ~x258 ;
  assign n494 = x2 & x258 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n492 & ~n495 ;
  assign n497 = ~n492 & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = n453 & n498 ;
  assign n500 = ~n453 & ~n498 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = ~n410 & n413 ;
  assign n503 = ~n414 & ~n502 ;
  assign n504 = n501 & n503 ;
  assign n505 = ~n414 & ~n504 ;
  assign n506 = n408 & ~n505 ;
  assign n507 = ~n433 & ~n451 ;
  assign n508 = ~n422 & ~n428 ;
  assign n509 = ~n507 & n508 ;
  assign n510 = n507 & ~n508 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = ~n443 & ~n449 ;
  assign n513 = n511 & n512 ;
  assign n514 = ~n511 & ~n512 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = ~n472 & ~n490 ;
  assign n517 = ~n461 & ~n467 ;
  assign n518 = ~n516 & n517 ;
  assign n519 = n516 & ~n517 ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = ~n482 & ~n488 ;
  assign n522 = n520 & n521 ;
  assign n523 = ~n520 & ~n521 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n496 & ~n499 ;
  assign n526 = n524 & ~n525 ;
  assign n527 = ~n524 & n525 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = n515 & n528 ;
  assign n530 = ~n515 & ~n528 ;
  assign n531 = ~n529 & ~n530 ;
  assign n532 = ~n408 & n505 ;
  assign n533 = ~n506 & ~n532 ;
  assign n534 = n531 & n533 ;
  assign n535 = ~n506 & ~n534 ;
  assign n536 = n406 & ~n535 ;
  assign n537 = ~n518 & ~n522 ;
  assign n538 = ~n526 & ~n529 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = n537 & n538 ;
  assign n541 = ~n539 & ~n540 ;
  assign n542 = ~n509 & ~n513 ;
  assign n543 = n541 & ~n542 ;
  assign n544 = ~n541 & n542 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~n406 & n535 ;
  assign n547 = ~n536 & ~n546 ;
  assign n548 = n545 & n547 ;
  assign n549 = ~n536 & ~n548 ;
  assign n550 = ~n404 & ~n549 ;
  assign n551 = n404 & n549 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = ~n539 & ~n543 ;
  assign n554 = n552 & ~n553 ;
  assign n555 = ~n552 & n553 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = ~n545 & ~n547 ;
  assign n558 = ~n548 & ~n557 ;
  assign n559 = ~n531 & ~n533 ;
  assign n560 = ~n534 & ~n559 ;
  assign n561 = ~n501 & ~n503 ;
  assign n562 = ~n504 & ~n561 ;
  assign n563 = ~x0 & ~x256 ;
  assign n564 = x0 & x256 ;
  assign n565 = ~n563 & ~n564 ;
  assign n566 = ~n562 & n565 ;
  assign n567 = ~n560 & n566 ;
  assign n568 = ~n558 & n567 ;
  assign n569 = ~n556 & n568 ;
  assign n570 = ~n550 & ~n554 ;
  assign n571 = n569 & n570 ;
  assign n572 = ~x254 & ~x286 ;
  assign n573 = x254 & x286 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = ~x253 & ~x285 ;
  assign n576 = x253 & x285 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = n574 & n577 ;
  assign n579 = ~n574 & ~n577 ;
  assign n580 = ~n578 & ~n579 ;
  assign n581 = ~x255 & ~x287 ;
  assign n582 = x255 & x287 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n580 & n583 ;
  assign n585 = ~n578 & ~n584 ;
  assign n586 = ~n580 & ~n583 ;
  assign n587 = ~n584 & ~n586 ;
  assign n588 = ~x249 & ~x281 ;
  assign n589 = x249 & x281 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = n587 & n590 ;
  assign n592 = ~x251 & ~x283 ;
  assign n593 = x251 & x283 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~x250 & ~x282 ;
  assign n596 = x250 & x282 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = ~n594 & ~n597 ;
  assign n599 = n594 & n597 ;
  assign n600 = ~n598 & ~n599 ;
  assign n601 = ~x252 & ~x284 ;
  assign n602 = x252 & x284 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = ~n600 & ~n603 ;
  assign n605 = n600 & n603 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = ~n587 & ~n590 ;
  assign n608 = ~n591 & ~n607 ;
  assign n609 = n606 & n608 ;
  assign n610 = ~n591 & ~n609 ;
  assign n611 = n585 & n610 ;
  assign n612 = ~n585 & ~n610 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = ~n599 & ~n605 ;
  assign n615 = n613 & n614 ;
  assign n616 = ~n611 & ~n615 ;
  assign n617 = ~n613 & ~n614 ;
  assign n618 = ~n615 & ~n617 ;
  assign n619 = ~n606 & ~n608 ;
  assign n620 = ~n609 & ~n619 ;
  assign n621 = ~x241 & ~x273 ;
  assign n622 = x241 & x273 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = n620 & n623 ;
  assign n625 = ~x247 & ~x279 ;
  assign n626 = x247 & x279 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~x246 & ~x278 ;
  assign n629 = x246 & x278 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = ~n627 & ~n630 ;
  assign n632 = n627 & n630 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = ~x248 & ~x280 ;
  assign n635 = x248 & x280 ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = ~n633 & ~n636 ;
  assign n638 = n633 & n636 ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = ~x242 & ~x274 ;
  assign n641 = x242 & x274 ;
  assign n642 = ~n640 & ~n641 ;
  assign n643 = ~n639 & ~n642 ;
  assign n644 = n639 & n642 ;
  assign n645 = ~n643 & ~n644 ;
  assign n646 = ~x244 & ~x276 ;
  assign n647 = x244 & x276 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = ~x243 & ~x275 ;
  assign n650 = x243 & x275 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = ~n648 & ~n651 ;
  assign n653 = n648 & n651 ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = ~x245 & ~x277 ;
  assign n656 = x245 & x277 ;
  assign n657 = ~n655 & ~n656 ;
  assign n658 = ~n654 & ~n657 ;
  assign n659 = n654 & n657 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = n645 & ~n660 ;
  assign n662 = ~n645 & n660 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = ~n620 & ~n623 ;
  assign n665 = ~n624 & ~n664 ;
  assign n666 = ~n663 & n665 ;
  assign n667 = ~n624 & ~n666 ;
  assign n668 = n618 & n667 ;
  assign n669 = ~n618 & ~n667 ;
  assign n670 = ~n643 & ~n661 ;
  assign n671 = ~n632 & ~n638 ;
  assign n672 = ~n670 & n671 ;
  assign n673 = n670 & ~n671 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~n653 & ~n659 ;
  assign n676 = n674 & n675 ;
  assign n677 = ~n674 & ~n675 ;
  assign n678 = ~n676 & ~n677 ;
  assign n679 = ~n669 & n678 ;
  assign n680 = ~n668 & ~n679 ;
  assign n681 = ~n616 & ~n680 ;
  assign n682 = n616 & n680 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = ~n672 & ~n676 ;
  assign n685 = n683 & ~n684 ;
  assign n686 = ~n681 & ~n685 ;
  assign n687 = ~n683 & n684 ;
  assign n688 = ~n685 & ~n687 ;
  assign n689 = n663 & ~n665 ;
  assign n690 = ~n666 & ~n689 ;
  assign n691 = ~x225 & ~x257 ;
  assign n692 = x225 & x257 ;
  assign n693 = ~n691 & ~n692 ;
  assign n694 = n690 & n693 ;
  assign n695 = ~x232 & ~x264 ;
  assign n696 = x232 & x264 ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = ~x231 & ~x263 ;
  assign n699 = x231 & x263 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~n697 & ~n700 ;
  assign n702 = n697 & n700 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~x233 & ~x265 ;
  assign n705 = x233 & x265 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n703 & ~n706 ;
  assign n708 = n703 & n706 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~x227 & ~x259 ;
  assign n711 = x227 & x259 ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = ~n709 & ~n712 ;
  assign n714 = n709 & n712 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~x229 & ~x261 ;
  assign n717 = x229 & x261 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~x228 & ~x260 ;
  assign n720 = x228 & x260 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~n718 & ~n721 ;
  assign n723 = n718 & n721 ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = ~x230 & ~x262 ;
  assign n726 = x230 & x262 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = ~n724 & ~n727 ;
  assign n729 = n724 & n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = n715 & ~n730 ;
  assign n732 = ~n715 & n730 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = ~x239 & ~x271 ;
  assign n735 = x239 & x271 ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = ~x238 & ~x270 ;
  assign n738 = x238 & x270 ;
  assign n739 = ~n737 & ~n738 ;
  assign n740 = ~n736 & ~n739 ;
  assign n741 = n736 & n739 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = ~x240 & ~x272 ;
  assign n744 = x240 & x272 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = ~n742 & ~n745 ;
  assign n747 = n742 & n745 ;
  assign n748 = ~n746 & ~n747 ;
  assign n749 = ~x234 & ~x266 ;
  assign n750 = x234 & x266 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~n748 & ~n751 ;
  assign n753 = n748 & n751 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~x236 & ~x268 ;
  assign n756 = x236 & x268 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = ~x235 & ~x267 ;
  assign n759 = x235 & x267 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = ~n757 & ~n760 ;
  assign n762 = n757 & n760 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~x237 & ~x269 ;
  assign n765 = x237 & x269 ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = ~n763 & ~n766 ;
  assign n768 = n763 & n766 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = n754 & ~n769 ;
  assign n771 = ~n754 & n769 ;
  assign n772 = ~n770 & ~n771 ;
  assign n773 = ~x226 & ~x258 ;
  assign n774 = x226 & x258 ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = n772 & ~n775 ;
  assign n777 = ~n772 & n775 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = n733 & n778 ;
  assign n780 = ~n733 & ~n778 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = ~n690 & ~n693 ;
  assign n783 = ~n694 & ~n782 ;
  assign n784 = ~n781 & n783 ;
  assign n785 = ~n694 & ~n784 ;
  assign n786 = ~n668 & ~n669 ;
  assign n787 = n678 & n786 ;
  assign n788 = ~n678 & ~n786 ;
  assign n789 = ~n787 & ~n788 ;
  assign n790 = ~n785 & ~n789 ;
  assign n791 = n785 & n789 ;
  assign n792 = ~n713 & ~n731 ;
  assign n793 = ~n702 & ~n708 ;
  assign n794 = ~n792 & n793 ;
  assign n795 = n792 & ~n793 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = ~n723 & ~n729 ;
  assign n798 = n796 & n797 ;
  assign n799 = ~n796 & ~n797 ;
  assign n800 = ~n798 & ~n799 ;
  assign n801 = ~n752 & ~n770 ;
  assign n802 = ~n741 & ~n747 ;
  assign n803 = ~n801 & n802 ;
  assign n804 = n801 & ~n802 ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = ~n762 & ~n768 ;
  assign n807 = n805 & n806 ;
  assign n808 = ~n805 & ~n806 ;
  assign n809 = ~n807 & ~n808 ;
  assign n810 = ~n776 & ~n779 ;
  assign n811 = n809 & ~n810 ;
  assign n812 = ~n809 & n810 ;
  assign n813 = ~n811 & ~n812 ;
  assign n814 = n800 & ~n813 ;
  assign n815 = ~n800 & n813 ;
  assign n816 = ~n814 & ~n815 ;
  assign n817 = ~n791 & n816 ;
  assign n818 = ~n790 & ~n817 ;
  assign n819 = ~n688 & ~n818 ;
  assign n820 = n688 & n818 ;
  assign n821 = ~n803 & ~n807 ;
  assign n822 = ~n812 & ~n815 ;
  assign n823 = ~n821 & n822 ;
  assign n824 = n821 & ~n822 ;
  assign n825 = ~n823 & ~n824 ;
  assign n826 = ~n794 & ~n798 ;
  assign n827 = n825 & ~n826 ;
  assign n828 = ~n825 & n826 ;
  assign n829 = ~n827 & ~n828 ;
  assign n830 = ~n820 & ~n829 ;
  assign n831 = ~n819 & ~n830 ;
  assign n832 = ~n686 & n831 ;
  assign n833 = n686 & ~n831 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = ~n823 & ~n827 ;
  assign n836 = n834 & ~n835 ;
  assign n837 = ~n832 & ~n836 ;
  assign n838 = ~n834 & n835 ;
  assign n839 = ~n836 & ~n838 ;
  assign n840 = n781 & ~n783 ;
  assign n841 = ~n784 & ~n840 ;
  assign n842 = ~x224 & ~x256 ;
  assign n843 = x224 & x256 ;
  assign n844 = ~n842 & ~n843 ;
  assign n845 = n841 & n844 ;
  assign n846 = ~n790 & ~n791 ;
  assign n847 = n816 & n846 ;
  assign n848 = ~n816 & ~n846 ;
  assign n849 = ~n847 & ~n848 ;
  assign n850 = n845 & n849 ;
  assign n851 = ~n819 & ~n820 ;
  assign n852 = ~n829 & n851 ;
  assign n853 = n829 & ~n851 ;
  assign n854 = ~n852 & ~n853 ;
  assign n855 = n850 & n854 ;
  assign n856 = ~n839 & n855 ;
  assign n857 = n837 & n856 ;
  assign n858 = ~x222 & ~x286 ;
  assign n859 = x222 & x286 ;
  assign n860 = ~n858 & ~n859 ;
  assign n861 = ~x221 & ~x285 ;
  assign n862 = x221 & x285 ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = n860 & n863 ;
  assign n865 = ~n860 & ~n863 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = ~x223 & ~x287 ;
  assign n868 = x223 & x287 ;
  assign n869 = ~n867 & ~n868 ;
  assign n870 = n866 & n869 ;
  assign n871 = ~n864 & ~n870 ;
  assign n872 = ~n866 & ~n869 ;
  assign n873 = ~n870 & ~n872 ;
  assign n874 = ~x217 & ~x281 ;
  assign n875 = x217 & x281 ;
  assign n876 = ~n874 & ~n875 ;
  assign n877 = n873 & n876 ;
  assign n878 = ~n873 & ~n876 ;
  assign n879 = ~x219 & ~x283 ;
  assign n880 = x219 & x283 ;
  assign n881 = ~n879 & ~n880 ;
  assign n882 = ~x218 & ~x282 ;
  assign n883 = x218 & x282 ;
  assign n884 = ~n882 & ~n883 ;
  assign n885 = ~n881 & ~n884 ;
  assign n886 = n881 & n884 ;
  assign n887 = ~n885 & ~n886 ;
  assign n888 = ~x220 & ~x284 ;
  assign n889 = x220 & x284 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = ~n887 & ~n890 ;
  assign n892 = n887 & n890 ;
  assign n893 = ~n891 & ~n892 ;
  assign n894 = ~n878 & n893 ;
  assign n895 = ~n877 & ~n894 ;
  assign n896 = n871 & n895 ;
  assign n897 = ~n871 & ~n895 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~n886 & ~n892 ;
  assign n900 = n898 & n899 ;
  assign n901 = ~n896 & ~n900 ;
  assign n902 = ~n898 & ~n899 ;
  assign n903 = ~n900 & ~n902 ;
  assign n904 = ~n877 & ~n878 ;
  assign n905 = ~n893 & n904 ;
  assign n906 = n893 & ~n904 ;
  assign n907 = ~n905 & ~n906 ;
  assign n908 = ~x209 & ~x273 ;
  assign n909 = x209 & x273 ;
  assign n910 = ~n908 & ~n909 ;
  assign n911 = ~n907 & n910 ;
  assign n912 = n907 & ~n910 ;
  assign n913 = ~x215 & ~x279 ;
  assign n914 = x215 & x279 ;
  assign n915 = ~n913 & ~n914 ;
  assign n916 = ~x214 & ~x278 ;
  assign n917 = x214 & x278 ;
  assign n918 = ~n916 & ~n917 ;
  assign n919 = ~n915 & ~n918 ;
  assign n920 = n915 & n918 ;
  assign n921 = ~n919 & ~n920 ;
  assign n922 = ~x216 & ~x280 ;
  assign n923 = x216 & x280 ;
  assign n924 = ~n922 & ~n923 ;
  assign n925 = ~n921 & ~n924 ;
  assign n926 = n921 & n924 ;
  assign n927 = ~n925 & ~n926 ;
  assign n928 = ~x210 & ~x274 ;
  assign n929 = x210 & x274 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = ~n927 & ~n930 ;
  assign n932 = n927 & n930 ;
  assign n933 = ~n931 & ~n932 ;
  assign n934 = ~x212 & ~x276 ;
  assign n935 = x212 & x276 ;
  assign n936 = ~n934 & ~n935 ;
  assign n937 = ~x211 & ~x275 ;
  assign n938 = x211 & x275 ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = ~n936 & ~n939 ;
  assign n941 = n936 & n939 ;
  assign n942 = ~n940 & ~n941 ;
  assign n943 = ~x213 & ~x277 ;
  assign n944 = x213 & x277 ;
  assign n945 = ~n943 & ~n944 ;
  assign n946 = ~n942 & ~n945 ;
  assign n947 = n942 & n945 ;
  assign n948 = ~n946 & ~n947 ;
  assign n949 = n933 & ~n948 ;
  assign n950 = ~n933 & n948 ;
  assign n951 = ~n949 & ~n950 ;
  assign n952 = ~n912 & ~n951 ;
  assign n953 = ~n911 & ~n952 ;
  assign n954 = n903 & n953 ;
  assign n955 = ~n903 & ~n953 ;
  assign n956 = ~n931 & ~n949 ;
  assign n957 = ~n920 & ~n926 ;
  assign n958 = ~n956 & n957 ;
  assign n959 = n956 & ~n957 ;
  assign n960 = ~n958 & ~n959 ;
  assign n961 = ~n941 & ~n947 ;
  assign n962 = n960 & n961 ;
  assign n963 = ~n960 & ~n961 ;
  assign n964 = ~n962 & ~n963 ;
  assign n965 = ~n955 & n964 ;
  assign n966 = ~n954 & ~n965 ;
  assign n967 = ~n901 & ~n966 ;
  assign n968 = n901 & n966 ;
  assign n969 = ~n967 & ~n968 ;
  assign n970 = ~n958 & ~n962 ;
  assign n971 = n969 & ~n970 ;
  assign n972 = ~n967 & ~n971 ;
  assign n973 = ~n969 & n970 ;
  assign n974 = ~n971 & ~n973 ;
  assign n975 = ~x193 & ~x257 ;
  assign n976 = x193 & x257 ;
  assign n977 = ~n975 & ~n976 ;
  assign n978 = ~n911 & ~n912 ;
  assign n979 = ~n951 & n978 ;
  assign n980 = n951 & ~n978 ;
  assign n981 = ~n979 & ~n980 ;
  assign n982 = ~n977 & ~n981 ;
  assign n983 = n977 & n981 ;
  assign n984 = ~x200 & ~x264 ;
  assign n985 = x200 & x264 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~x199 & ~x263 ;
  assign n988 = x199 & x263 ;
  assign n989 = ~n987 & ~n988 ;
  assign n990 = ~n986 & ~n989 ;
  assign n991 = n986 & n989 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = ~x201 & ~x265 ;
  assign n994 = x201 & x265 ;
  assign n995 = ~n993 & ~n994 ;
  assign n996 = ~n992 & ~n995 ;
  assign n997 = n992 & n995 ;
  assign n998 = ~n996 & ~n997 ;
  assign n999 = ~x195 & ~x259 ;
  assign n1000 = x195 & x259 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1002 = ~n998 & ~n1001 ;
  assign n1003 = n998 & n1001 ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = ~x197 & ~x261 ;
  assign n1006 = x197 & x261 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = ~x196 & ~x260 ;
  assign n1009 = x196 & x260 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = ~n1007 & ~n1010 ;
  assign n1012 = n1007 & n1010 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = ~x198 & ~x262 ;
  assign n1015 = x198 & x262 ;
  assign n1016 = ~n1014 & ~n1015 ;
  assign n1017 = ~n1013 & ~n1016 ;
  assign n1018 = n1013 & n1016 ;
  assign n1019 = ~n1017 & ~n1018 ;
  assign n1020 = n1004 & ~n1019 ;
  assign n1021 = ~n1004 & n1019 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = ~x207 & ~x271 ;
  assign n1024 = x207 & x271 ;
  assign n1025 = ~n1023 & ~n1024 ;
  assign n1026 = ~x206 & ~x270 ;
  assign n1027 = x206 & x270 ;
  assign n1028 = ~n1026 & ~n1027 ;
  assign n1029 = ~n1025 & ~n1028 ;
  assign n1030 = n1025 & n1028 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = ~x208 & ~x272 ;
  assign n1033 = x208 & x272 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = ~n1031 & ~n1034 ;
  assign n1036 = n1031 & n1034 ;
  assign n1037 = ~n1035 & ~n1036 ;
  assign n1038 = ~x202 & ~x266 ;
  assign n1039 = x202 & x266 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1041 = ~n1037 & ~n1040 ;
  assign n1042 = n1037 & n1040 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = ~x204 & ~x268 ;
  assign n1045 = x204 & x268 ;
  assign n1046 = ~n1044 & ~n1045 ;
  assign n1047 = ~x203 & ~x267 ;
  assign n1048 = x203 & x267 ;
  assign n1049 = ~n1047 & ~n1048 ;
  assign n1050 = ~n1046 & ~n1049 ;
  assign n1051 = n1046 & n1049 ;
  assign n1052 = ~n1050 & ~n1051 ;
  assign n1053 = ~x205 & ~x269 ;
  assign n1054 = x205 & x269 ;
  assign n1055 = ~n1053 & ~n1054 ;
  assign n1056 = ~n1052 & ~n1055 ;
  assign n1057 = n1052 & n1055 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = n1043 & ~n1058 ;
  assign n1060 = ~n1043 & n1058 ;
  assign n1061 = ~n1059 & ~n1060 ;
  assign n1062 = ~x194 & ~x258 ;
  assign n1063 = x194 & x258 ;
  assign n1064 = ~n1062 & ~n1063 ;
  assign n1065 = n1061 & ~n1064 ;
  assign n1066 = ~n1061 & n1064 ;
  assign n1067 = ~n1065 & ~n1066 ;
  assign n1068 = n1022 & n1067 ;
  assign n1069 = ~n1022 & ~n1067 ;
  assign n1070 = ~n1068 & ~n1069 ;
  assign n1071 = ~n983 & n1070 ;
  assign n1072 = ~n982 & ~n1071 ;
  assign n1073 = ~n954 & ~n955 ;
  assign n1074 = ~n964 & n1073 ;
  assign n1075 = n964 & ~n1073 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1077 = n1072 & n1076 ;
  assign n1078 = ~n1072 & ~n1076 ;
  assign n1079 = ~n1002 & ~n1020 ;
  assign n1080 = ~n991 & ~n997 ;
  assign n1081 = ~n1079 & n1080 ;
  assign n1082 = n1079 & ~n1080 ;
  assign n1083 = ~n1081 & ~n1082 ;
  assign n1084 = ~n1012 & ~n1018 ;
  assign n1085 = n1083 & n1084 ;
  assign n1086 = ~n1083 & ~n1084 ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1088 = ~n1041 & ~n1059 ;
  assign n1089 = ~n1030 & ~n1036 ;
  assign n1090 = ~n1088 & n1089 ;
  assign n1091 = n1088 & ~n1089 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = ~n1051 & ~n1057 ;
  assign n1094 = n1092 & n1093 ;
  assign n1095 = ~n1092 & ~n1093 ;
  assign n1096 = ~n1094 & ~n1095 ;
  assign n1097 = ~n1065 & ~n1068 ;
  assign n1098 = n1096 & ~n1097 ;
  assign n1099 = ~n1096 & n1097 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = n1087 & n1100 ;
  assign n1102 = ~n1087 & ~n1100 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = ~n1078 & ~n1103 ;
  assign n1105 = ~n1077 & ~n1104 ;
  assign n1106 = ~n974 & ~n1105 ;
  assign n1107 = n974 & n1105 ;
  assign n1108 = ~n1087 & ~n1098 ;
  assign n1109 = ~n1099 & ~n1108 ;
  assign n1110 = ~n1090 & ~n1094 ;
  assign n1111 = n1109 & ~n1110 ;
  assign n1112 = ~n1109 & n1110 ;
  assign n1113 = ~n1111 & ~n1112 ;
  assign n1114 = ~n1081 & ~n1085 ;
  assign n1115 = n1113 & ~n1114 ;
  assign n1116 = ~n1113 & n1114 ;
  assign n1117 = ~n1115 & ~n1116 ;
  assign n1118 = ~n1107 & ~n1117 ;
  assign n1119 = ~n1106 & ~n1118 ;
  assign n1120 = ~n972 & n1119 ;
  assign n1121 = n972 & ~n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~n1111 & ~n1115 ;
  assign n1124 = n1122 & ~n1123 ;
  assign n1125 = ~n1120 & ~n1124 ;
  assign n1126 = ~n1122 & n1123 ;
  assign n1127 = ~n1124 & ~n1126 ;
  assign n1128 = ~x192 & ~x256 ;
  assign n1129 = x192 & x256 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1131 = ~n982 & ~n983 ;
  assign n1132 = n1070 & n1131 ;
  assign n1133 = ~n1070 & ~n1131 ;
  assign n1134 = ~n1132 & ~n1133 ;
  assign n1135 = n1130 & ~n1134 ;
  assign n1136 = ~n1077 & ~n1078 ;
  assign n1137 = ~n1103 & n1136 ;
  assign n1138 = n1103 & ~n1136 ;
  assign n1139 = ~n1137 & ~n1138 ;
  assign n1140 = n1135 & n1139 ;
  assign n1141 = ~n1106 & ~n1107 ;
  assign n1142 = ~n1117 & n1141 ;
  assign n1143 = n1117 & ~n1141 ;
  assign n1144 = ~n1142 & ~n1143 ;
  assign n1145 = n1140 & n1144 ;
  assign n1146 = ~n1127 & n1145 ;
  assign n1147 = n1125 & n1146 ;
  assign n1148 = n857 & n1147 ;
  assign n1149 = ~x190 & ~x286 ;
  assign n1150 = x190 & x286 ;
  assign n1151 = ~n1149 & ~n1150 ;
  assign n1152 = ~x189 & ~x285 ;
  assign n1153 = x189 & x285 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = n1151 & n1154 ;
  assign n1156 = ~n1151 & ~n1154 ;
  assign n1157 = ~n1155 & ~n1156 ;
  assign n1158 = ~x191 & ~x287 ;
  assign n1159 = x191 & x287 ;
  assign n1160 = ~n1158 & ~n1159 ;
  assign n1161 = ~n1157 & ~n1160 ;
  assign n1162 = n1157 & n1160 ;
  assign n1163 = ~n1161 & ~n1162 ;
  assign n1164 = ~x185 & ~x281 ;
  assign n1165 = x185 & x281 ;
  assign n1166 = ~n1164 & ~n1165 ;
  assign n1167 = ~n1163 & ~n1166 ;
  assign n1168 = n1163 & n1166 ;
  assign n1169 = ~n1167 & ~n1168 ;
  assign n1170 = ~x187 & ~x283 ;
  assign n1171 = x187 & x283 ;
  assign n1172 = ~n1170 & ~n1171 ;
  assign n1173 = ~x186 & ~x282 ;
  assign n1174 = x186 & x282 ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1176 = ~n1172 & ~n1175 ;
  assign n1177 = n1172 & n1175 ;
  assign n1178 = ~n1176 & ~n1177 ;
  assign n1179 = ~x188 & ~x284 ;
  assign n1180 = x188 & x284 ;
  assign n1181 = ~n1179 & ~n1180 ;
  assign n1182 = ~n1178 & ~n1181 ;
  assign n1183 = n1178 & n1181 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = n1169 & ~n1184 ;
  assign n1186 = ~n1167 & ~n1185 ;
  assign n1187 = ~n1155 & ~n1162 ;
  assign n1188 = ~n1186 & n1187 ;
  assign n1189 = n1186 & ~n1187 ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = ~n1177 & ~n1183 ;
  assign n1192 = n1190 & n1191 ;
  assign n1193 = ~n1188 & ~n1192 ;
  assign n1194 = ~n1190 & ~n1191 ;
  assign n1195 = ~n1192 & ~n1194 ;
  assign n1196 = ~n1169 & n1184 ;
  assign n1197 = ~n1185 & ~n1196 ;
  assign n1198 = ~x177 & ~x273 ;
  assign n1199 = x177 & x273 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1201 = n1197 & ~n1200 ;
  assign n1202 = ~x183 & ~x279 ;
  assign n1203 = x183 & x279 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1205 = ~x182 & ~x278 ;
  assign n1206 = x182 & x278 ;
  assign n1207 = ~n1205 & ~n1206 ;
  assign n1208 = ~n1204 & ~n1207 ;
  assign n1209 = n1204 & n1207 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = ~x184 & ~x280 ;
  assign n1212 = x184 & x280 ;
  assign n1213 = ~n1211 & ~n1212 ;
  assign n1214 = ~n1210 & ~n1213 ;
  assign n1215 = n1210 & n1213 ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = ~x178 & ~x274 ;
  assign n1218 = x178 & x274 ;
  assign n1219 = ~n1217 & ~n1218 ;
  assign n1220 = ~n1216 & ~n1219 ;
  assign n1221 = n1216 & n1219 ;
  assign n1222 = ~n1220 & ~n1221 ;
  assign n1223 = ~x180 & ~x276 ;
  assign n1224 = x180 & x276 ;
  assign n1225 = ~n1223 & ~n1224 ;
  assign n1226 = ~x179 & ~x275 ;
  assign n1227 = x179 & x275 ;
  assign n1228 = ~n1226 & ~n1227 ;
  assign n1229 = ~n1225 & ~n1228 ;
  assign n1230 = n1225 & n1228 ;
  assign n1231 = ~n1229 & ~n1230 ;
  assign n1232 = ~x181 & ~x277 ;
  assign n1233 = x181 & x277 ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = ~n1231 & ~n1234 ;
  assign n1236 = n1231 & n1234 ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = n1222 & ~n1237 ;
  assign n1239 = ~n1222 & n1237 ;
  assign n1240 = ~n1238 & ~n1239 ;
  assign n1241 = ~n1197 & n1200 ;
  assign n1242 = ~n1201 & ~n1241 ;
  assign n1243 = n1240 & n1242 ;
  assign n1244 = ~n1201 & ~n1243 ;
  assign n1245 = n1195 & ~n1244 ;
  assign n1246 = ~n1220 & ~n1238 ;
  assign n1247 = ~n1209 & ~n1215 ;
  assign n1248 = ~n1246 & n1247 ;
  assign n1249 = n1246 & ~n1247 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = ~n1230 & ~n1236 ;
  assign n1252 = n1250 & n1251 ;
  assign n1253 = ~n1250 & ~n1251 ;
  assign n1254 = ~n1252 & ~n1253 ;
  assign n1255 = ~n1195 & n1244 ;
  assign n1256 = ~n1245 & ~n1255 ;
  assign n1257 = n1254 & n1256 ;
  assign n1258 = ~n1245 & ~n1257 ;
  assign n1259 = ~n1193 & ~n1258 ;
  assign n1260 = n1193 & n1258 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = ~n1248 & ~n1252 ;
  assign n1263 = n1261 & ~n1262 ;
  assign n1264 = ~n1259 & ~n1263 ;
  assign n1265 = ~n1261 & n1262 ;
  assign n1266 = ~n1263 & ~n1265 ;
  assign n1267 = ~n1254 & ~n1256 ;
  assign n1268 = ~n1257 & ~n1267 ;
  assign n1269 = ~n1240 & ~n1242 ;
  assign n1270 = ~n1243 & ~n1269 ;
  assign n1271 = ~x161 & ~x257 ;
  assign n1272 = x161 & x257 ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = n1270 & ~n1273 ;
  assign n1275 = ~x168 & ~x264 ;
  assign n1276 = x168 & x264 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = ~x167 & ~x263 ;
  assign n1279 = x167 & x263 ;
  assign n1280 = ~n1278 & ~n1279 ;
  assign n1281 = ~n1277 & ~n1280 ;
  assign n1282 = n1277 & n1280 ;
  assign n1283 = ~n1281 & ~n1282 ;
  assign n1284 = ~x169 & ~x265 ;
  assign n1285 = x169 & x265 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = ~n1283 & ~n1286 ;
  assign n1288 = n1283 & n1286 ;
  assign n1289 = ~n1287 & ~n1288 ;
  assign n1290 = ~x163 & ~x259 ;
  assign n1291 = x163 & x259 ;
  assign n1292 = ~n1290 & ~n1291 ;
  assign n1293 = ~n1289 & ~n1292 ;
  assign n1294 = n1289 & n1292 ;
  assign n1295 = ~n1293 & ~n1294 ;
  assign n1296 = ~x165 & ~x261 ;
  assign n1297 = x165 & x261 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = ~x164 & ~x260 ;
  assign n1300 = x164 & x260 ;
  assign n1301 = ~n1299 & ~n1300 ;
  assign n1302 = ~n1298 & ~n1301 ;
  assign n1303 = n1298 & n1301 ;
  assign n1304 = ~n1302 & ~n1303 ;
  assign n1305 = ~x166 & ~x262 ;
  assign n1306 = x166 & x262 ;
  assign n1307 = ~n1305 & ~n1306 ;
  assign n1308 = ~n1304 & ~n1307 ;
  assign n1309 = n1304 & n1307 ;
  assign n1310 = ~n1308 & ~n1309 ;
  assign n1311 = n1295 & ~n1310 ;
  assign n1312 = ~n1295 & n1310 ;
  assign n1313 = ~n1311 & ~n1312 ;
  assign n1314 = ~x175 & ~x271 ;
  assign n1315 = x175 & x271 ;
  assign n1316 = ~n1314 & ~n1315 ;
  assign n1317 = ~x174 & ~x270 ;
  assign n1318 = x174 & x270 ;
  assign n1319 = ~n1317 & ~n1318 ;
  assign n1320 = ~n1316 & ~n1319 ;
  assign n1321 = n1316 & n1319 ;
  assign n1322 = ~n1320 & ~n1321 ;
  assign n1323 = ~x176 & ~x272 ;
  assign n1324 = x176 & x272 ;
  assign n1325 = ~n1323 & ~n1324 ;
  assign n1326 = ~n1322 & ~n1325 ;
  assign n1327 = n1322 & n1325 ;
  assign n1328 = ~n1326 & ~n1327 ;
  assign n1329 = ~x170 & ~x266 ;
  assign n1330 = x170 & x266 ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = ~n1328 & ~n1331 ;
  assign n1333 = n1328 & n1331 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = ~x172 & ~x268 ;
  assign n1336 = x172 & x268 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = ~x171 & ~x267 ;
  assign n1339 = x171 & x267 ;
  assign n1340 = ~n1338 & ~n1339 ;
  assign n1341 = ~n1337 & ~n1340 ;
  assign n1342 = n1337 & n1340 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = ~x173 & ~x269 ;
  assign n1345 = x173 & x269 ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = ~n1343 & ~n1346 ;
  assign n1348 = n1343 & n1346 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = n1334 & ~n1349 ;
  assign n1351 = ~n1334 & n1349 ;
  assign n1352 = ~n1350 & ~n1351 ;
  assign n1353 = ~x162 & ~x258 ;
  assign n1354 = x162 & x258 ;
  assign n1355 = ~n1353 & ~n1354 ;
  assign n1356 = n1352 & ~n1355 ;
  assign n1357 = ~n1352 & n1355 ;
  assign n1358 = ~n1356 & ~n1357 ;
  assign n1359 = n1313 & n1358 ;
  assign n1360 = ~n1313 & ~n1358 ;
  assign n1361 = ~n1359 & ~n1360 ;
  assign n1362 = ~n1270 & n1273 ;
  assign n1363 = ~n1274 & ~n1362 ;
  assign n1364 = n1361 & n1363 ;
  assign n1365 = ~n1274 & ~n1364 ;
  assign n1366 = n1268 & ~n1365 ;
  assign n1367 = ~n1293 & ~n1311 ;
  assign n1368 = ~n1282 & ~n1288 ;
  assign n1369 = ~n1367 & n1368 ;
  assign n1370 = n1367 & ~n1368 ;
  assign n1371 = ~n1369 & ~n1370 ;
  assign n1372 = ~n1303 & ~n1309 ;
  assign n1373 = n1371 & n1372 ;
  assign n1374 = ~n1371 & ~n1372 ;
  assign n1375 = ~n1373 & ~n1374 ;
  assign n1376 = ~n1332 & ~n1350 ;
  assign n1377 = ~n1321 & ~n1327 ;
  assign n1378 = ~n1376 & n1377 ;
  assign n1379 = n1376 & ~n1377 ;
  assign n1380 = ~n1378 & ~n1379 ;
  assign n1381 = ~n1342 & ~n1348 ;
  assign n1382 = n1380 & n1381 ;
  assign n1383 = ~n1380 & ~n1381 ;
  assign n1384 = ~n1382 & ~n1383 ;
  assign n1385 = ~n1356 & ~n1359 ;
  assign n1386 = n1384 & ~n1385 ;
  assign n1387 = ~n1384 & n1385 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = n1375 & n1388 ;
  assign n1390 = ~n1375 & ~n1388 ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1392 = ~n1268 & n1365 ;
  assign n1393 = ~n1366 & ~n1392 ;
  assign n1394 = n1391 & n1393 ;
  assign n1395 = ~n1366 & ~n1394 ;
  assign n1396 = n1266 & ~n1395 ;
  assign n1397 = ~n1378 & ~n1382 ;
  assign n1398 = ~n1386 & ~n1389 ;
  assign n1399 = ~n1397 & ~n1398 ;
  assign n1400 = n1397 & n1398 ;
  assign n1401 = ~n1399 & ~n1400 ;
  assign n1402 = ~n1369 & ~n1373 ;
  assign n1403 = n1401 & ~n1402 ;
  assign n1404 = ~n1401 & n1402 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~n1266 & n1395 ;
  assign n1407 = ~n1396 & ~n1406 ;
  assign n1408 = n1405 & n1407 ;
  assign n1409 = ~n1396 & ~n1408 ;
  assign n1410 = ~n1264 & ~n1409 ;
  assign n1411 = n1264 & n1409 ;
  assign n1412 = ~n1410 & ~n1411 ;
  assign n1413 = ~n1399 & ~n1403 ;
  assign n1414 = n1412 & ~n1413 ;
  assign n1415 = ~n1410 & ~n1414 ;
  assign n1416 = ~n1412 & n1413 ;
  assign n1417 = ~n1414 & ~n1416 ;
  assign n1418 = ~n1405 & ~n1407 ;
  assign n1419 = ~n1408 & ~n1418 ;
  assign n1420 = ~n1391 & ~n1393 ;
  assign n1421 = ~n1394 & ~n1420 ;
  assign n1422 = ~n1361 & ~n1363 ;
  assign n1423 = ~n1364 & ~n1422 ;
  assign n1424 = ~x160 & ~x256 ;
  assign n1425 = x160 & x256 ;
  assign n1426 = ~n1424 & ~n1425 ;
  assign n1427 = ~n1423 & n1426 ;
  assign n1428 = ~n1421 & n1427 ;
  assign n1429 = ~n1419 & n1428 ;
  assign n1430 = ~n1417 & n1429 ;
  assign n1431 = n1415 & n1430 ;
  assign n1432 = n1148 & n1431 ;
  assign n1433 = ~x158 & ~x286 ;
  assign n1434 = x158 & x286 ;
  assign n1435 = ~n1433 & ~n1434 ;
  assign n1436 = ~x157 & ~x285 ;
  assign n1437 = x157 & x285 ;
  assign n1438 = ~n1436 & ~n1437 ;
  assign n1439 = n1435 & n1438 ;
  assign n1440 = ~n1435 & ~n1438 ;
  assign n1441 = ~n1439 & ~n1440 ;
  assign n1442 = ~x159 & ~x287 ;
  assign n1443 = x159 & x287 ;
  assign n1444 = ~n1442 & ~n1443 ;
  assign n1445 = ~n1441 & ~n1444 ;
  assign n1446 = n1441 & n1444 ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1448 = ~x153 & ~x281 ;
  assign n1449 = x153 & x281 ;
  assign n1450 = ~n1448 & ~n1449 ;
  assign n1451 = ~n1447 & ~n1450 ;
  assign n1452 = n1447 & n1450 ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = ~x155 & ~x283 ;
  assign n1455 = x155 & x283 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = ~x154 & ~x282 ;
  assign n1458 = x154 & x282 ;
  assign n1459 = ~n1457 & ~n1458 ;
  assign n1460 = ~n1456 & ~n1459 ;
  assign n1461 = n1456 & n1459 ;
  assign n1462 = ~n1460 & ~n1461 ;
  assign n1463 = ~x156 & ~x284 ;
  assign n1464 = x156 & x284 ;
  assign n1465 = ~n1463 & ~n1464 ;
  assign n1466 = ~n1462 & ~n1465 ;
  assign n1467 = n1462 & n1465 ;
  assign n1468 = ~n1466 & ~n1467 ;
  assign n1469 = n1453 & ~n1468 ;
  assign n1470 = ~n1451 & ~n1469 ;
  assign n1471 = ~n1439 & ~n1446 ;
  assign n1472 = ~n1470 & n1471 ;
  assign n1473 = n1470 & ~n1471 ;
  assign n1474 = ~n1472 & ~n1473 ;
  assign n1475 = ~n1461 & ~n1467 ;
  assign n1476 = n1474 & n1475 ;
  assign n1477 = ~n1472 & ~n1476 ;
  assign n1478 = ~n1474 & ~n1475 ;
  assign n1479 = ~n1476 & ~n1478 ;
  assign n1480 = ~n1453 & n1468 ;
  assign n1481 = ~n1469 & ~n1480 ;
  assign n1482 = ~x145 & ~x273 ;
  assign n1483 = x145 & x273 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = n1481 & ~n1484 ;
  assign n1486 = ~x151 & ~x279 ;
  assign n1487 = x151 & x279 ;
  assign n1488 = ~n1486 & ~n1487 ;
  assign n1489 = ~x150 & ~x278 ;
  assign n1490 = x150 & x278 ;
  assign n1491 = ~n1489 & ~n1490 ;
  assign n1492 = ~n1488 & ~n1491 ;
  assign n1493 = n1488 & n1491 ;
  assign n1494 = ~n1492 & ~n1493 ;
  assign n1495 = ~x152 & ~x280 ;
  assign n1496 = x152 & x280 ;
  assign n1497 = ~n1495 & ~n1496 ;
  assign n1498 = ~n1494 & ~n1497 ;
  assign n1499 = n1494 & n1497 ;
  assign n1500 = ~n1498 & ~n1499 ;
  assign n1501 = ~x146 & ~x274 ;
  assign n1502 = x146 & x274 ;
  assign n1503 = ~n1501 & ~n1502 ;
  assign n1504 = ~n1500 & ~n1503 ;
  assign n1505 = n1500 & n1503 ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = ~x148 & ~x276 ;
  assign n1508 = x148 & x276 ;
  assign n1509 = ~n1507 & ~n1508 ;
  assign n1510 = ~x147 & ~x275 ;
  assign n1511 = x147 & x275 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = ~n1509 & ~n1512 ;
  assign n1514 = n1509 & n1512 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = ~x149 & ~x277 ;
  assign n1517 = x149 & x277 ;
  assign n1518 = ~n1516 & ~n1517 ;
  assign n1519 = ~n1515 & ~n1518 ;
  assign n1520 = n1515 & n1518 ;
  assign n1521 = ~n1519 & ~n1520 ;
  assign n1522 = n1506 & ~n1521 ;
  assign n1523 = ~n1506 & n1521 ;
  assign n1524 = ~n1522 & ~n1523 ;
  assign n1525 = ~n1481 & n1484 ;
  assign n1526 = ~n1485 & ~n1525 ;
  assign n1527 = n1524 & n1526 ;
  assign n1528 = ~n1485 & ~n1527 ;
  assign n1529 = n1479 & ~n1528 ;
  assign n1530 = ~n1504 & ~n1522 ;
  assign n1531 = ~n1493 & ~n1499 ;
  assign n1532 = ~n1530 & n1531 ;
  assign n1533 = n1530 & ~n1531 ;
  assign n1534 = ~n1532 & ~n1533 ;
  assign n1535 = ~n1514 & ~n1520 ;
  assign n1536 = n1534 & n1535 ;
  assign n1537 = ~n1534 & ~n1535 ;
  assign n1538 = ~n1536 & ~n1537 ;
  assign n1539 = ~n1479 & n1528 ;
  assign n1540 = ~n1529 & ~n1539 ;
  assign n1541 = n1538 & n1540 ;
  assign n1542 = ~n1529 & ~n1541 ;
  assign n1543 = ~n1477 & ~n1542 ;
  assign n1544 = n1477 & n1542 ;
  assign n1545 = ~n1543 & ~n1544 ;
  assign n1546 = ~n1532 & ~n1536 ;
  assign n1547 = n1545 & ~n1546 ;
  assign n1548 = ~n1543 & ~n1547 ;
  assign n1549 = ~n1545 & n1546 ;
  assign n1550 = ~n1547 & ~n1549 ;
  assign n1551 = ~n1538 & ~n1540 ;
  assign n1552 = ~n1541 & ~n1551 ;
  assign n1553 = ~n1524 & ~n1526 ;
  assign n1554 = ~n1527 & ~n1553 ;
  assign n1555 = ~x129 & ~x257 ;
  assign n1556 = x129 & x257 ;
  assign n1557 = ~n1555 & ~n1556 ;
  assign n1558 = n1554 & ~n1557 ;
  assign n1559 = ~x136 & ~x264 ;
  assign n1560 = x136 & x264 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~x135 & ~x263 ;
  assign n1563 = x135 & x263 ;
  assign n1564 = ~n1562 & ~n1563 ;
  assign n1565 = ~n1561 & ~n1564 ;
  assign n1566 = n1561 & n1564 ;
  assign n1567 = ~n1565 & ~n1566 ;
  assign n1568 = ~x137 & ~x265 ;
  assign n1569 = x137 & x265 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1571 = ~n1567 & ~n1570 ;
  assign n1572 = n1567 & n1570 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = ~x131 & ~x259 ;
  assign n1575 = x131 & x259 ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = ~n1573 & ~n1576 ;
  assign n1578 = n1573 & n1576 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = ~x133 & ~x261 ;
  assign n1581 = x133 & x261 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = ~x132 & ~x260 ;
  assign n1584 = x132 & x260 ;
  assign n1585 = ~n1583 & ~n1584 ;
  assign n1586 = ~n1582 & ~n1585 ;
  assign n1587 = n1582 & n1585 ;
  assign n1588 = ~n1586 & ~n1587 ;
  assign n1589 = ~x134 & ~x262 ;
  assign n1590 = x134 & x262 ;
  assign n1591 = ~n1589 & ~n1590 ;
  assign n1592 = ~n1588 & ~n1591 ;
  assign n1593 = n1588 & n1591 ;
  assign n1594 = ~n1592 & ~n1593 ;
  assign n1595 = n1579 & ~n1594 ;
  assign n1596 = ~n1579 & n1594 ;
  assign n1597 = ~n1595 & ~n1596 ;
  assign n1598 = ~x143 & ~x271 ;
  assign n1599 = x143 & x271 ;
  assign n1600 = ~n1598 & ~n1599 ;
  assign n1601 = ~x142 & ~x270 ;
  assign n1602 = x142 & x270 ;
  assign n1603 = ~n1601 & ~n1602 ;
  assign n1604 = ~n1600 & ~n1603 ;
  assign n1605 = n1600 & n1603 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1607 = ~x144 & ~x272 ;
  assign n1608 = x144 & x272 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = ~n1606 & ~n1609 ;
  assign n1611 = n1606 & n1609 ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1613 = ~x138 & ~x266 ;
  assign n1614 = x138 & x266 ;
  assign n1615 = ~n1613 & ~n1614 ;
  assign n1616 = ~n1612 & ~n1615 ;
  assign n1617 = n1612 & n1615 ;
  assign n1618 = ~n1616 & ~n1617 ;
  assign n1619 = ~x140 & ~x268 ;
  assign n1620 = x140 & x268 ;
  assign n1621 = ~n1619 & ~n1620 ;
  assign n1622 = ~x139 & ~x267 ;
  assign n1623 = x139 & x267 ;
  assign n1624 = ~n1622 & ~n1623 ;
  assign n1625 = ~n1621 & ~n1624 ;
  assign n1626 = n1621 & n1624 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = ~x141 & ~x269 ;
  assign n1629 = x141 & x269 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = ~n1627 & ~n1630 ;
  assign n1632 = n1627 & n1630 ;
  assign n1633 = ~n1631 & ~n1632 ;
  assign n1634 = n1618 & ~n1633 ;
  assign n1635 = ~n1618 & n1633 ;
  assign n1636 = ~n1634 & ~n1635 ;
  assign n1637 = ~x130 & ~x258 ;
  assign n1638 = x130 & x258 ;
  assign n1639 = ~n1637 & ~n1638 ;
  assign n1640 = n1636 & ~n1639 ;
  assign n1641 = ~n1636 & n1639 ;
  assign n1642 = ~n1640 & ~n1641 ;
  assign n1643 = n1597 & n1642 ;
  assign n1644 = ~n1597 & ~n1642 ;
  assign n1645 = ~n1643 & ~n1644 ;
  assign n1646 = ~n1554 & n1557 ;
  assign n1647 = ~n1558 & ~n1646 ;
  assign n1648 = n1645 & n1647 ;
  assign n1649 = ~n1558 & ~n1648 ;
  assign n1650 = n1552 & ~n1649 ;
  assign n1651 = ~n1577 & ~n1595 ;
  assign n1652 = ~n1566 & ~n1572 ;
  assign n1653 = ~n1651 & n1652 ;
  assign n1654 = n1651 & ~n1652 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = ~n1587 & ~n1593 ;
  assign n1657 = n1655 & n1656 ;
  assign n1658 = ~n1655 & ~n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = ~n1616 & ~n1634 ;
  assign n1661 = ~n1605 & ~n1611 ;
  assign n1662 = ~n1660 & n1661 ;
  assign n1663 = n1660 & ~n1661 ;
  assign n1664 = ~n1662 & ~n1663 ;
  assign n1665 = ~n1626 & ~n1632 ;
  assign n1666 = n1664 & n1665 ;
  assign n1667 = ~n1664 & ~n1665 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1669 = ~n1640 & ~n1643 ;
  assign n1670 = n1668 & ~n1669 ;
  assign n1671 = ~n1668 & n1669 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = n1659 & n1672 ;
  assign n1674 = ~n1659 & ~n1672 ;
  assign n1675 = ~n1673 & ~n1674 ;
  assign n1676 = ~n1552 & n1649 ;
  assign n1677 = ~n1650 & ~n1676 ;
  assign n1678 = n1675 & n1677 ;
  assign n1679 = ~n1650 & ~n1678 ;
  assign n1680 = n1550 & ~n1679 ;
  assign n1681 = ~n1662 & ~n1666 ;
  assign n1682 = ~n1670 & ~n1673 ;
  assign n1683 = ~n1681 & ~n1682 ;
  assign n1684 = n1681 & n1682 ;
  assign n1685 = ~n1683 & ~n1684 ;
  assign n1686 = ~n1653 & ~n1657 ;
  assign n1687 = n1685 & ~n1686 ;
  assign n1688 = ~n1685 & n1686 ;
  assign n1689 = ~n1687 & ~n1688 ;
  assign n1690 = ~n1550 & n1679 ;
  assign n1691 = ~n1680 & ~n1690 ;
  assign n1692 = n1689 & n1691 ;
  assign n1693 = ~n1680 & ~n1692 ;
  assign n1694 = ~n1548 & ~n1693 ;
  assign n1695 = n1548 & n1693 ;
  assign n1696 = ~n1694 & ~n1695 ;
  assign n1697 = ~n1683 & ~n1687 ;
  assign n1698 = n1696 & ~n1697 ;
  assign n1699 = ~n1694 & ~n1698 ;
  assign n1700 = ~n1696 & n1697 ;
  assign n1701 = ~n1698 & ~n1700 ;
  assign n1702 = ~n1689 & ~n1691 ;
  assign n1703 = ~n1692 & ~n1702 ;
  assign n1704 = ~n1675 & ~n1677 ;
  assign n1705 = ~n1678 & ~n1704 ;
  assign n1706 = ~n1645 & ~n1647 ;
  assign n1707 = ~n1648 & ~n1706 ;
  assign n1708 = ~x128 & ~x256 ;
  assign n1709 = x128 & x256 ;
  assign n1710 = ~n1708 & ~n1709 ;
  assign n1711 = ~n1707 & n1710 ;
  assign n1712 = ~n1705 & n1711 ;
  assign n1713 = ~n1703 & n1712 ;
  assign n1714 = ~n1701 & n1713 ;
  assign n1715 = n1699 & n1714 ;
  assign n1716 = n1432 & n1715 ;
  assign n1717 = ~x126 & ~x286 ;
  assign n1718 = x126 & x286 ;
  assign n1719 = ~n1717 & ~n1718 ;
  assign n1720 = ~x125 & ~x285 ;
  assign n1721 = x125 & x285 ;
  assign n1722 = ~n1720 & ~n1721 ;
  assign n1723 = n1719 & n1722 ;
  assign n1724 = ~n1719 & ~n1722 ;
  assign n1725 = ~n1723 & ~n1724 ;
  assign n1726 = ~x127 & ~x287 ;
  assign n1727 = x127 & x287 ;
  assign n1728 = ~n1726 & ~n1727 ;
  assign n1729 = ~n1725 & ~n1728 ;
  assign n1730 = n1725 & n1728 ;
  assign n1731 = ~n1729 & ~n1730 ;
  assign n1732 = ~x121 & ~x281 ;
  assign n1733 = x121 & x281 ;
  assign n1734 = ~n1732 & ~n1733 ;
  assign n1735 = ~n1731 & ~n1734 ;
  assign n1736 = n1731 & n1734 ;
  assign n1737 = ~n1735 & ~n1736 ;
  assign n1738 = ~x123 & ~x283 ;
  assign n1739 = x123 & x283 ;
  assign n1740 = ~n1738 & ~n1739 ;
  assign n1741 = ~x122 & ~x282 ;
  assign n1742 = x122 & x282 ;
  assign n1743 = ~n1741 & ~n1742 ;
  assign n1744 = ~n1740 & ~n1743 ;
  assign n1745 = n1740 & n1743 ;
  assign n1746 = ~n1744 & ~n1745 ;
  assign n1747 = ~x124 & ~x284 ;
  assign n1748 = x124 & x284 ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = ~n1746 & ~n1749 ;
  assign n1751 = n1746 & n1749 ;
  assign n1752 = ~n1750 & ~n1751 ;
  assign n1753 = n1737 & ~n1752 ;
  assign n1754 = ~n1735 & ~n1753 ;
  assign n1755 = ~n1723 & ~n1730 ;
  assign n1756 = ~n1754 & n1755 ;
  assign n1757 = n1754 & ~n1755 ;
  assign n1758 = ~n1756 & ~n1757 ;
  assign n1759 = ~n1745 & ~n1751 ;
  assign n1760 = n1758 & n1759 ;
  assign n1761 = ~n1756 & ~n1760 ;
  assign n1762 = ~n1758 & ~n1759 ;
  assign n1763 = ~n1760 & ~n1762 ;
  assign n1764 = ~n1737 & n1752 ;
  assign n1765 = ~n1753 & ~n1764 ;
  assign n1766 = ~x113 & ~x273 ;
  assign n1767 = x113 & x273 ;
  assign n1768 = ~n1766 & ~n1767 ;
  assign n1769 = n1765 & ~n1768 ;
  assign n1770 = ~x119 & ~x279 ;
  assign n1771 = x119 & x279 ;
  assign n1772 = ~n1770 & ~n1771 ;
  assign n1773 = ~x118 & ~x278 ;
  assign n1774 = x118 & x278 ;
  assign n1775 = ~n1773 & ~n1774 ;
  assign n1776 = ~n1772 & ~n1775 ;
  assign n1777 = n1772 & n1775 ;
  assign n1778 = ~n1776 & ~n1777 ;
  assign n1779 = ~x120 & ~x280 ;
  assign n1780 = x120 & x280 ;
  assign n1781 = ~n1779 & ~n1780 ;
  assign n1782 = ~n1778 & ~n1781 ;
  assign n1783 = n1778 & n1781 ;
  assign n1784 = ~n1782 & ~n1783 ;
  assign n1785 = ~x114 & ~x274 ;
  assign n1786 = x114 & x274 ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1788 = ~n1784 & ~n1787 ;
  assign n1789 = n1784 & n1787 ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1791 = ~x116 & ~x276 ;
  assign n1792 = x116 & x276 ;
  assign n1793 = ~n1791 & ~n1792 ;
  assign n1794 = ~x115 & ~x275 ;
  assign n1795 = x115 & x275 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = ~n1793 & ~n1796 ;
  assign n1798 = n1793 & n1796 ;
  assign n1799 = ~n1797 & ~n1798 ;
  assign n1800 = ~x117 & ~x277 ;
  assign n1801 = x117 & x277 ;
  assign n1802 = ~n1800 & ~n1801 ;
  assign n1803 = ~n1799 & ~n1802 ;
  assign n1804 = n1799 & n1802 ;
  assign n1805 = ~n1803 & ~n1804 ;
  assign n1806 = n1790 & ~n1805 ;
  assign n1807 = ~n1790 & n1805 ;
  assign n1808 = ~n1806 & ~n1807 ;
  assign n1809 = ~n1765 & n1768 ;
  assign n1810 = ~n1769 & ~n1809 ;
  assign n1811 = n1808 & n1810 ;
  assign n1812 = ~n1769 & ~n1811 ;
  assign n1813 = n1763 & ~n1812 ;
  assign n1814 = ~n1788 & ~n1806 ;
  assign n1815 = ~n1777 & ~n1783 ;
  assign n1816 = ~n1814 & n1815 ;
  assign n1817 = n1814 & ~n1815 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = ~n1798 & ~n1804 ;
  assign n1820 = n1818 & n1819 ;
  assign n1821 = ~n1818 & ~n1819 ;
  assign n1822 = ~n1820 & ~n1821 ;
  assign n1823 = ~n1763 & n1812 ;
  assign n1824 = ~n1813 & ~n1823 ;
  assign n1825 = n1822 & n1824 ;
  assign n1826 = ~n1813 & ~n1825 ;
  assign n1827 = ~n1761 & ~n1826 ;
  assign n1828 = n1761 & n1826 ;
  assign n1829 = ~n1827 & ~n1828 ;
  assign n1830 = ~n1816 & ~n1820 ;
  assign n1831 = n1829 & ~n1830 ;
  assign n1832 = ~n1827 & ~n1831 ;
  assign n1833 = ~n1829 & n1830 ;
  assign n1834 = ~n1831 & ~n1833 ;
  assign n1835 = ~n1822 & ~n1824 ;
  assign n1836 = ~n1825 & ~n1835 ;
  assign n1837 = ~n1808 & ~n1810 ;
  assign n1838 = ~n1811 & ~n1837 ;
  assign n1839 = ~x97 & ~x257 ;
  assign n1840 = x97 & x257 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = n1838 & ~n1841 ;
  assign n1843 = ~x104 & ~x264 ;
  assign n1844 = x104 & x264 ;
  assign n1845 = ~n1843 & ~n1844 ;
  assign n1846 = ~x103 & ~x263 ;
  assign n1847 = x103 & x263 ;
  assign n1848 = ~n1846 & ~n1847 ;
  assign n1849 = ~n1845 & ~n1848 ;
  assign n1850 = n1845 & n1848 ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = ~x105 & ~x265 ;
  assign n1853 = x105 & x265 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = ~n1851 & ~n1854 ;
  assign n1856 = n1851 & n1854 ;
  assign n1857 = ~n1855 & ~n1856 ;
  assign n1858 = ~x99 & ~x259 ;
  assign n1859 = x99 & x259 ;
  assign n1860 = ~n1858 & ~n1859 ;
  assign n1861 = ~n1857 & ~n1860 ;
  assign n1862 = n1857 & n1860 ;
  assign n1863 = ~n1861 & ~n1862 ;
  assign n1864 = ~x101 & ~x261 ;
  assign n1865 = x101 & x261 ;
  assign n1866 = ~n1864 & ~n1865 ;
  assign n1867 = ~x100 & ~x260 ;
  assign n1868 = x100 & x260 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1870 = ~n1866 & ~n1869 ;
  assign n1871 = n1866 & n1869 ;
  assign n1872 = ~n1870 & ~n1871 ;
  assign n1873 = ~x102 & ~x262 ;
  assign n1874 = x102 & x262 ;
  assign n1875 = ~n1873 & ~n1874 ;
  assign n1876 = ~n1872 & ~n1875 ;
  assign n1877 = n1872 & n1875 ;
  assign n1878 = ~n1876 & ~n1877 ;
  assign n1879 = n1863 & ~n1878 ;
  assign n1880 = ~n1863 & n1878 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = ~x111 & ~x271 ;
  assign n1883 = x111 & x271 ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1885 = ~x110 & ~x270 ;
  assign n1886 = x110 & x270 ;
  assign n1887 = ~n1885 & ~n1886 ;
  assign n1888 = ~n1884 & ~n1887 ;
  assign n1889 = n1884 & n1887 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = ~x112 & ~x272 ;
  assign n1892 = x112 & x272 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = ~n1890 & ~n1893 ;
  assign n1895 = n1890 & n1893 ;
  assign n1896 = ~n1894 & ~n1895 ;
  assign n1897 = ~x106 & ~x266 ;
  assign n1898 = x106 & x266 ;
  assign n1899 = ~n1897 & ~n1898 ;
  assign n1900 = ~n1896 & ~n1899 ;
  assign n1901 = n1896 & n1899 ;
  assign n1902 = ~n1900 & ~n1901 ;
  assign n1903 = ~x108 & ~x268 ;
  assign n1904 = x108 & x268 ;
  assign n1905 = ~n1903 & ~n1904 ;
  assign n1906 = ~x107 & ~x267 ;
  assign n1907 = x107 & x267 ;
  assign n1908 = ~n1906 & ~n1907 ;
  assign n1909 = ~n1905 & ~n1908 ;
  assign n1910 = n1905 & n1908 ;
  assign n1911 = ~n1909 & ~n1910 ;
  assign n1912 = ~x109 & ~x269 ;
  assign n1913 = x109 & x269 ;
  assign n1914 = ~n1912 & ~n1913 ;
  assign n1915 = ~n1911 & ~n1914 ;
  assign n1916 = n1911 & n1914 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = n1902 & ~n1917 ;
  assign n1919 = ~n1902 & n1917 ;
  assign n1920 = ~n1918 & ~n1919 ;
  assign n1921 = ~x98 & ~x258 ;
  assign n1922 = x98 & x258 ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1924 = n1920 & ~n1923 ;
  assign n1925 = ~n1920 & n1923 ;
  assign n1926 = ~n1924 & ~n1925 ;
  assign n1927 = n1881 & n1926 ;
  assign n1928 = ~n1881 & ~n1926 ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1930 = ~n1838 & n1841 ;
  assign n1931 = ~n1842 & ~n1930 ;
  assign n1932 = n1929 & n1931 ;
  assign n1933 = ~n1842 & ~n1932 ;
  assign n1934 = n1836 & ~n1933 ;
  assign n1935 = ~n1861 & ~n1879 ;
  assign n1936 = ~n1850 & ~n1856 ;
  assign n1937 = ~n1935 & n1936 ;
  assign n1938 = n1935 & ~n1936 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = ~n1871 & ~n1877 ;
  assign n1941 = n1939 & n1940 ;
  assign n1942 = ~n1939 & ~n1940 ;
  assign n1943 = ~n1941 & ~n1942 ;
  assign n1944 = ~n1900 & ~n1918 ;
  assign n1945 = ~n1889 & ~n1895 ;
  assign n1946 = ~n1944 & n1945 ;
  assign n1947 = n1944 & ~n1945 ;
  assign n1948 = ~n1946 & ~n1947 ;
  assign n1949 = ~n1910 & ~n1916 ;
  assign n1950 = n1948 & n1949 ;
  assign n1951 = ~n1948 & ~n1949 ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1953 = ~n1924 & ~n1927 ;
  assign n1954 = n1952 & ~n1953 ;
  assign n1955 = ~n1952 & n1953 ;
  assign n1956 = ~n1954 & ~n1955 ;
  assign n1957 = n1943 & n1956 ;
  assign n1958 = ~n1943 & ~n1956 ;
  assign n1959 = ~n1957 & ~n1958 ;
  assign n1960 = ~n1836 & n1933 ;
  assign n1961 = ~n1934 & ~n1960 ;
  assign n1962 = n1959 & n1961 ;
  assign n1963 = ~n1934 & ~n1962 ;
  assign n1964 = n1834 & ~n1963 ;
  assign n1965 = ~n1946 & ~n1950 ;
  assign n1966 = ~n1954 & ~n1957 ;
  assign n1967 = ~n1965 & ~n1966 ;
  assign n1968 = n1965 & n1966 ;
  assign n1969 = ~n1967 & ~n1968 ;
  assign n1970 = ~n1937 & ~n1941 ;
  assign n1971 = n1969 & ~n1970 ;
  assign n1972 = ~n1969 & n1970 ;
  assign n1973 = ~n1971 & ~n1972 ;
  assign n1974 = ~n1834 & n1963 ;
  assign n1975 = ~n1964 & ~n1974 ;
  assign n1976 = n1973 & n1975 ;
  assign n1977 = ~n1964 & ~n1976 ;
  assign n1978 = ~n1832 & ~n1977 ;
  assign n1979 = n1832 & n1977 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = ~n1967 & ~n1971 ;
  assign n1982 = n1980 & ~n1981 ;
  assign n1983 = ~n1978 & ~n1982 ;
  assign n1984 = ~n1980 & n1981 ;
  assign n1985 = ~n1982 & ~n1984 ;
  assign n1986 = ~n1973 & ~n1975 ;
  assign n1987 = ~n1976 & ~n1986 ;
  assign n1988 = ~n1959 & ~n1961 ;
  assign n1989 = ~n1962 & ~n1988 ;
  assign n1990 = ~n1929 & ~n1931 ;
  assign n1991 = ~n1932 & ~n1990 ;
  assign n1992 = ~x96 & ~x256 ;
  assign n1993 = x96 & x256 ;
  assign n1994 = ~n1992 & ~n1993 ;
  assign n1995 = ~n1991 & n1994 ;
  assign n1996 = ~n1989 & n1995 ;
  assign n1997 = ~n1987 & n1996 ;
  assign n1998 = ~n1985 & n1997 ;
  assign n1999 = n1983 & n1998 ;
  assign n2000 = n1716 & n1999 ;
  assign n2001 = ~x94 & ~x286 ;
  assign n2002 = x94 & x286 ;
  assign n2003 = ~n2001 & ~n2002 ;
  assign n2004 = ~x93 & ~x285 ;
  assign n2005 = x93 & x285 ;
  assign n2006 = ~n2004 & ~n2005 ;
  assign n2007 = n2003 & n2006 ;
  assign n2008 = ~n2003 & ~n2006 ;
  assign n2009 = ~n2007 & ~n2008 ;
  assign n2010 = ~x95 & ~x287 ;
  assign n2011 = x95 & x287 ;
  assign n2012 = ~n2010 & ~n2011 ;
  assign n2013 = ~n2009 & ~n2012 ;
  assign n2014 = n2009 & n2012 ;
  assign n2015 = ~n2013 & ~n2014 ;
  assign n2016 = ~x89 & ~x281 ;
  assign n2017 = x89 & x281 ;
  assign n2018 = ~n2016 & ~n2017 ;
  assign n2019 = ~n2015 & ~n2018 ;
  assign n2020 = n2015 & n2018 ;
  assign n2021 = ~n2019 & ~n2020 ;
  assign n2022 = ~x91 & ~x283 ;
  assign n2023 = x91 & x283 ;
  assign n2024 = ~n2022 & ~n2023 ;
  assign n2025 = ~x90 & ~x282 ;
  assign n2026 = x90 & x282 ;
  assign n2027 = ~n2025 & ~n2026 ;
  assign n2028 = ~n2024 & ~n2027 ;
  assign n2029 = n2024 & n2027 ;
  assign n2030 = ~n2028 & ~n2029 ;
  assign n2031 = ~x92 & ~x284 ;
  assign n2032 = x92 & x284 ;
  assign n2033 = ~n2031 & ~n2032 ;
  assign n2034 = ~n2030 & ~n2033 ;
  assign n2035 = n2030 & n2033 ;
  assign n2036 = ~n2034 & ~n2035 ;
  assign n2037 = n2021 & ~n2036 ;
  assign n2038 = ~n2019 & ~n2037 ;
  assign n2039 = ~n2007 & ~n2014 ;
  assign n2040 = ~n2038 & n2039 ;
  assign n2041 = n2038 & ~n2039 ;
  assign n2042 = ~n2040 & ~n2041 ;
  assign n2043 = ~n2029 & ~n2035 ;
  assign n2044 = n2042 & n2043 ;
  assign n2045 = ~n2040 & ~n2044 ;
  assign n2046 = ~n2042 & ~n2043 ;
  assign n2047 = ~n2044 & ~n2046 ;
  assign n2048 = ~n2021 & n2036 ;
  assign n2049 = ~n2037 & ~n2048 ;
  assign n2050 = ~x81 & ~x273 ;
  assign n2051 = x81 & x273 ;
  assign n2052 = ~n2050 & ~n2051 ;
  assign n2053 = n2049 & ~n2052 ;
  assign n2054 = ~x87 & ~x279 ;
  assign n2055 = x87 & x279 ;
  assign n2056 = ~n2054 & ~n2055 ;
  assign n2057 = ~x86 & ~x278 ;
  assign n2058 = x86 & x278 ;
  assign n2059 = ~n2057 & ~n2058 ;
  assign n2060 = ~n2056 & ~n2059 ;
  assign n2061 = n2056 & n2059 ;
  assign n2062 = ~n2060 & ~n2061 ;
  assign n2063 = ~x88 & ~x280 ;
  assign n2064 = x88 & x280 ;
  assign n2065 = ~n2063 & ~n2064 ;
  assign n2066 = ~n2062 & ~n2065 ;
  assign n2067 = n2062 & n2065 ;
  assign n2068 = ~n2066 & ~n2067 ;
  assign n2069 = ~x82 & ~x274 ;
  assign n2070 = x82 & x274 ;
  assign n2071 = ~n2069 & ~n2070 ;
  assign n2072 = ~n2068 & ~n2071 ;
  assign n2073 = n2068 & n2071 ;
  assign n2074 = ~n2072 & ~n2073 ;
  assign n2075 = ~x84 & ~x276 ;
  assign n2076 = x84 & x276 ;
  assign n2077 = ~n2075 & ~n2076 ;
  assign n2078 = ~x83 & ~x275 ;
  assign n2079 = x83 & x275 ;
  assign n2080 = ~n2078 & ~n2079 ;
  assign n2081 = ~n2077 & ~n2080 ;
  assign n2082 = n2077 & n2080 ;
  assign n2083 = ~n2081 & ~n2082 ;
  assign n2084 = ~x85 & ~x277 ;
  assign n2085 = x85 & x277 ;
  assign n2086 = ~n2084 & ~n2085 ;
  assign n2087 = ~n2083 & ~n2086 ;
  assign n2088 = n2083 & n2086 ;
  assign n2089 = ~n2087 & ~n2088 ;
  assign n2090 = n2074 & ~n2089 ;
  assign n2091 = ~n2074 & n2089 ;
  assign n2092 = ~n2090 & ~n2091 ;
  assign n2093 = ~n2049 & n2052 ;
  assign n2094 = ~n2053 & ~n2093 ;
  assign n2095 = n2092 & n2094 ;
  assign n2096 = ~n2053 & ~n2095 ;
  assign n2097 = n2047 & ~n2096 ;
  assign n2098 = ~n2072 & ~n2090 ;
  assign n2099 = ~n2061 & ~n2067 ;
  assign n2100 = ~n2098 & n2099 ;
  assign n2101 = n2098 & ~n2099 ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = ~n2082 & ~n2088 ;
  assign n2104 = n2102 & n2103 ;
  assign n2105 = ~n2102 & ~n2103 ;
  assign n2106 = ~n2104 & ~n2105 ;
  assign n2107 = ~n2047 & n2096 ;
  assign n2108 = ~n2097 & ~n2107 ;
  assign n2109 = n2106 & n2108 ;
  assign n2110 = ~n2097 & ~n2109 ;
  assign n2111 = ~n2045 & ~n2110 ;
  assign n2112 = n2045 & n2110 ;
  assign n2113 = ~n2111 & ~n2112 ;
  assign n2114 = ~n2100 & ~n2104 ;
  assign n2115 = n2113 & ~n2114 ;
  assign n2116 = ~n2111 & ~n2115 ;
  assign n2117 = ~n2113 & n2114 ;
  assign n2118 = ~n2115 & ~n2117 ;
  assign n2119 = ~n2106 & ~n2108 ;
  assign n2120 = ~n2109 & ~n2119 ;
  assign n2121 = ~n2092 & ~n2094 ;
  assign n2122 = ~n2095 & ~n2121 ;
  assign n2123 = ~x65 & ~x257 ;
  assign n2124 = x65 & x257 ;
  assign n2125 = ~n2123 & ~n2124 ;
  assign n2126 = n2122 & ~n2125 ;
  assign n2127 = ~x72 & ~x264 ;
  assign n2128 = x72 & x264 ;
  assign n2129 = ~n2127 & ~n2128 ;
  assign n2130 = ~x71 & ~x263 ;
  assign n2131 = x71 & x263 ;
  assign n2132 = ~n2130 & ~n2131 ;
  assign n2133 = ~n2129 & ~n2132 ;
  assign n2134 = n2129 & n2132 ;
  assign n2135 = ~n2133 & ~n2134 ;
  assign n2136 = ~x73 & ~x265 ;
  assign n2137 = x73 & x265 ;
  assign n2138 = ~n2136 & ~n2137 ;
  assign n2139 = ~n2135 & ~n2138 ;
  assign n2140 = n2135 & n2138 ;
  assign n2141 = ~n2139 & ~n2140 ;
  assign n2142 = ~x67 & ~x259 ;
  assign n2143 = x67 & x259 ;
  assign n2144 = ~n2142 & ~n2143 ;
  assign n2145 = ~n2141 & ~n2144 ;
  assign n2146 = n2141 & n2144 ;
  assign n2147 = ~n2145 & ~n2146 ;
  assign n2148 = ~x69 & ~x261 ;
  assign n2149 = x69 & x261 ;
  assign n2150 = ~n2148 & ~n2149 ;
  assign n2151 = ~x68 & ~x260 ;
  assign n2152 = x68 & x260 ;
  assign n2153 = ~n2151 & ~n2152 ;
  assign n2154 = ~n2150 & ~n2153 ;
  assign n2155 = n2150 & n2153 ;
  assign n2156 = ~n2154 & ~n2155 ;
  assign n2157 = ~x70 & ~x262 ;
  assign n2158 = x70 & x262 ;
  assign n2159 = ~n2157 & ~n2158 ;
  assign n2160 = ~n2156 & ~n2159 ;
  assign n2161 = n2156 & n2159 ;
  assign n2162 = ~n2160 & ~n2161 ;
  assign n2163 = n2147 & ~n2162 ;
  assign n2164 = ~n2147 & n2162 ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2166 = ~x79 & ~x271 ;
  assign n2167 = x79 & x271 ;
  assign n2168 = ~n2166 & ~n2167 ;
  assign n2169 = ~x78 & ~x270 ;
  assign n2170 = x78 & x270 ;
  assign n2171 = ~n2169 & ~n2170 ;
  assign n2172 = ~n2168 & ~n2171 ;
  assign n2173 = n2168 & n2171 ;
  assign n2174 = ~n2172 & ~n2173 ;
  assign n2175 = ~x80 & ~x272 ;
  assign n2176 = x80 & x272 ;
  assign n2177 = ~n2175 & ~n2176 ;
  assign n2178 = ~n2174 & ~n2177 ;
  assign n2179 = n2174 & n2177 ;
  assign n2180 = ~n2178 & ~n2179 ;
  assign n2181 = ~x74 & ~x266 ;
  assign n2182 = x74 & x266 ;
  assign n2183 = ~n2181 & ~n2182 ;
  assign n2184 = ~n2180 & ~n2183 ;
  assign n2185 = n2180 & n2183 ;
  assign n2186 = ~n2184 & ~n2185 ;
  assign n2187 = ~x76 & ~x268 ;
  assign n2188 = x76 & x268 ;
  assign n2189 = ~n2187 & ~n2188 ;
  assign n2190 = ~x75 & ~x267 ;
  assign n2191 = x75 & x267 ;
  assign n2192 = ~n2190 & ~n2191 ;
  assign n2193 = ~n2189 & ~n2192 ;
  assign n2194 = n2189 & n2192 ;
  assign n2195 = ~n2193 & ~n2194 ;
  assign n2196 = ~x77 & ~x269 ;
  assign n2197 = x77 & x269 ;
  assign n2198 = ~n2196 & ~n2197 ;
  assign n2199 = ~n2195 & ~n2198 ;
  assign n2200 = n2195 & n2198 ;
  assign n2201 = ~n2199 & ~n2200 ;
  assign n2202 = n2186 & ~n2201 ;
  assign n2203 = ~n2186 & n2201 ;
  assign n2204 = ~n2202 & ~n2203 ;
  assign n2205 = ~x66 & ~x258 ;
  assign n2206 = x66 & x258 ;
  assign n2207 = ~n2205 & ~n2206 ;
  assign n2208 = n2204 & ~n2207 ;
  assign n2209 = ~n2204 & n2207 ;
  assign n2210 = ~n2208 & ~n2209 ;
  assign n2211 = n2165 & n2210 ;
  assign n2212 = ~n2165 & ~n2210 ;
  assign n2213 = ~n2211 & ~n2212 ;
  assign n2214 = ~n2122 & n2125 ;
  assign n2215 = ~n2126 & ~n2214 ;
  assign n2216 = n2213 & n2215 ;
  assign n2217 = ~n2126 & ~n2216 ;
  assign n2218 = n2120 & ~n2217 ;
  assign n2219 = ~n2145 & ~n2163 ;
  assign n2220 = ~n2134 & ~n2140 ;
  assign n2221 = ~n2219 & n2220 ;
  assign n2222 = n2219 & ~n2220 ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = ~n2155 & ~n2161 ;
  assign n2225 = n2223 & n2224 ;
  assign n2226 = ~n2223 & ~n2224 ;
  assign n2227 = ~n2225 & ~n2226 ;
  assign n2228 = ~n2184 & ~n2202 ;
  assign n2229 = ~n2173 & ~n2179 ;
  assign n2230 = ~n2228 & n2229 ;
  assign n2231 = n2228 & ~n2229 ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = ~n2194 & ~n2200 ;
  assign n2234 = n2232 & n2233 ;
  assign n2235 = ~n2232 & ~n2233 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = ~n2208 & ~n2211 ;
  assign n2238 = n2236 & ~n2237 ;
  assign n2239 = ~n2236 & n2237 ;
  assign n2240 = ~n2238 & ~n2239 ;
  assign n2241 = n2227 & n2240 ;
  assign n2242 = ~n2227 & ~n2240 ;
  assign n2243 = ~n2241 & ~n2242 ;
  assign n2244 = ~n2120 & n2217 ;
  assign n2245 = ~n2218 & ~n2244 ;
  assign n2246 = n2243 & n2245 ;
  assign n2247 = ~n2218 & ~n2246 ;
  assign n2248 = n2118 & ~n2247 ;
  assign n2249 = ~n2230 & ~n2234 ;
  assign n2250 = ~n2238 & ~n2241 ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = n2249 & n2250 ;
  assign n2253 = ~n2251 & ~n2252 ;
  assign n2254 = ~n2221 & ~n2225 ;
  assign n2255 = n2253 & ~n2254 ;
  assign n2256 = ~n2253 & n2254 ;
  assign n2257 = ~n2255 & ~n2256 ;
  assign n2258 = ~n2118 & n2247 ;
  assign n2259 = ~n2248 & ~n2258 ;
  assign n2260 = n2257 & n2259 ;
  assign n2261 = ~n2248 & ~n2260 ;
  assign n2262 = ~n2116 & ~n2261 ;
  assign n2263 = n2116 & n2261 ;
  assign n2264 = ~n2262 & ~n2263 ;
  assign n2265 = ~n2251 & ~n2255 ;
  assign n2266 = n2264 & ~n2265 ;
  assign n2267 = ~n2262 & ~n2266 ;
  assign n2268 = ~n2264 & n2265 ;
  assign n2269 = ~n2266 & ~n2268 ;
  assign n2270 = ~n2257 & ~n2259 ;
  assign n2271 = ~n2260 & ~n2270 ;
  assign n2272 = ~n2213 & ~n2215 ;
  assign n2273 = ~n2216 & ~n2272 ;
  assign n2274 = ~x64 & ~x256 ;
  assign n2275 = x64 & x256 ;
  assign n2276 = ~n2274 & ~n2275 ;
  assign n2277 = ~n2273 & n2276 ;
  assign n2278 = ~n2243 & ~n2245 ;
  assign n2279 = ~n2246 & ~n2278 ;
  assign n2280 = n2277 & ~n2279 ;
  assign n2281 = ~n2271 & n2280 ;
  assign n2282 = ~n2269 & n2281 ;
  assign n2283 = n2267 & n2282 ;
  assign n2284 = n2000 & n2283 ;
  assign n2285 = ~x62 & ~x286 ;
  assign n2286 = x62 & x286 ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = ~x61 & ~x285 ;
  assign n2289 = x61 & x285 ;
  assign n2290 = ~n2288 & ~n2289 ;
  assign n2291 = ~n2287 & ~n2290 ;
  assign n2292 = n2287 & n2290 ;
  assign n2293 = ~n2291 & ~n2292 ;
  assign n2294 = ~x63 & ~x287 ;
  assign n2295 = x63 & x287 ;
  assign n2296 = ~n2294 & ~n2295 ;
  assign n2297 = ~n2293 & ~n2296 ;
  assign n2298 = n2293 & n2296 ;
  assign n2299 = ~n2297 & ~n2298 ;
  assign n2300 = ~x57 & ~x281 ;
  assign n2301 = x57 & x281 ;
  assign n2302 = ~n2300 & ~n2301 ;
  assign n2303 = ~n2299 & ~n2302 ;
  assign n2304 = n2299 & n2302 ;
  assign n2305 = ~n2303 & ~n2304 ;
  assign n2306 = ~x59 & ~x283 ;
  assign n2307 = x59 & x283 ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = ~x58 & ~x282 ;
  assign n2310 = x58 & x282 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = ~n2308 & ~n2311 ;
  assign n2313 = n2308 & n2311 ;
  assign n2314 = ~n2312 & ~n2313 ;
  assign n2315 = ~x60 & ~x284 ;
  assign n2316 = x60 & x284 ;
  assign n2317 = ~n2315 & ~n2316 ;
  assign n2318 = ~n2314 & ~n2317 ;
  assign n2319 = n2314 & n2317 ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = n2305 & ~n2320 ;
  assign n2322 = ~n2303 & ~n2321 ;
  assign n2323 = ~n2292 & ~n2298 ;
  assign n2324 = ~n2322 & n2323 ;
  assign n2325 = n2322 & ~n2323 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = ~n2313 & ~n2319 ;
  assign n2328 = n2326 & n2327 ;
  assign n2329 = ~n2324 & ~n2328 ;
  assign n2330 = ~n2326 & ~n2327 ;
  assign n2331 = ~n2328 & ~n2330 ;
  assign n2332 = ~n2305 & n2320 ;
  assign n2333 = ~n2321 & ~n2332 ;
  assign n2334 = ~x49 & ~x273 ;
  assign n2335 = x49 & x273 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = n2333 & ~n2336 ;
  assign n2338 = ~x55 & ~x279 ;
  assign n2339 = x55 & x279 ;
  assign n2340 = ~n2338 & ~n2339 ;
  assign n2341 = ~x54 & ~x278 ;
  assign n2342 = x54 & x278 ;
  assign n2343 = ~n2341 & ~n2342 ;
  assign n2344 = ~n2340 & ~n2343 ;
  assign n2345 = n2340 & n2343 ;
  assign n2346 = ~n2344 & ~n2345 ;
  assign n2347 = ~x56 & ~x280 ;
  assign n2348 = x56 & x280 ;
  assign n2349 = ~n2347 & ~n2348 ;
  assign n2350 = ~n2346 & ~n2349 ;
  assign n2351 = n2346 & n2349 ;
  assign n2352 = ~n2350 & ~n2351 ;
  assign n2353 = ~x50 & ~x274 ;
  assign n2354 = x50 & x274 ;
  assign n2355 = ~n2353 & ~n2354 ;
  assign n2356 = ~n2352 & ~n2355 ;
  assign n2357 = n2352 & n2355 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = ~x52 & ~x276 ;
  assign n2360 = x52 & x276 ;
  assign n2361 = ~n2359 & ~n2360 ;
  assign n2362 = ~x51 & ~x275 ;
  assign n2363 = x51 & x275 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = ~n2361 & ~n2364 ;
  assign n2366 = n2361 & n2364 ;
  assign n2367 = ~n2365 & ~n2366 ;
  assign n2368 = ~x53 & ~x277 ;
  assign n2369 = x53 & x277 ;
  assign n2370 = ~n2368 & ~n2369 ;
  assign n2371 = ~n2367 & ~n2370 ;
  assign n2372 = n2367 & n2370 ;
  assign n2373 = ~n2371 & ~n2372 ;
  assign n2374 = n2358 & ~n2373 ;
  assign n2375 = ~n2358 & n2373 ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2377 = ~n2333 & n2336 ;
  assign n2378 = ~n2337 & ~n2377 ;
  assign n2379 = n2376 & n2378 ;
  assign n2380 = ~n2337 & ~n2379 ;
  assign n2381 = n2331 & ~n2380 ;
  assign n2382 = ~n2356 & ~n2374 ;
  assign n2383 = ~n2345 & ~n2351 ;
  assign n2384 = ~n2382 & n2383 ;
  assign n2385 = n2382 & ~n2383 ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2387 = ~n2366 & ~n2372 ;
  assign n2388 = n2386 & n2387 ;
  assign n2389 = ~n2386 & ~n2387 ;
  assign n2390 = ~n2388 & ~n2389 ;
  assign n2391 = ~n2331 & n2380 ;
  assign n2392 = ~n2381 & ~n2391 ;
  assign n2393 = n2390 & n2392 ;
  assign n2394 = ~n2381 & ~n2393 ;
  assign n2395 = ~n2329 & ~n2394 ;
  assign n2396 = n2329 & n2394 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = ~n2384 & ~n2388 ;
  assign n2399 = n2397 & ~n2398 ;
  assign n2400 = ~n2395 & ~n2399 ;
  assign n2401 = ~n2397 & n2398 ;
  assign n2402 = ~n2399 & ~n2401 ;
  assign n2403 = ~n2390 & ~n2392 ;
  assign n2404 = ~n2393 & ~n2403 ;
  assign n2405 = ~n2376 & ~n2378 ;
  assign n2406 = ~n2379 & ~n2405 ;
  assign n2407 = ~x33 & ~x257 ;
  assign n2408 = x33 & x257 ;
  assign n2409 = ~n2407 & ~n2408 ;
  assign n2410 = n2406 & ~n2409 ;
  assign n2411 = ~x40 & ~x264 ;
  assign n2412 = x40 & x264 ;
  assign n2413 = ~n2411 & ~n2412 ;
  assign n2414 = ~x39 & ~x263 ;
  assign n2415 = x39 & x263 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = ~n2413 & ~n2416 ;
  assign n2418 = n2413 & n2416 ;
  assign n2419 = ~n2417 & ~n2418 ;
  assign n2420 = ~x41 & ~x265 ;
  assign n2421 = x41 & x265 ;
  assign n2422 = ~n2420 & ~n2421 ;
  assign n2423 = ~n2419 & ~n2422 ;
  assign n2424 = n2419 & n2422 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = ~x35 & ~x259 ;
  assign n2427 = x35 & x259 ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign n2429 = ~n2425 & ~n2428 ;
  assign n2430 = n2425 & n2428 ;
  assign n2431 = ~n2429 & ~n2430 ;
  assign n2432 = ~x37 & ~x261 ;
  assign n2433 = x37 & x261 ;
  assign n2434 = ~n2432 & ~n2433 ;
  assign n2435 = ~x36 & ~x260 ;
  assign n2436 = x36 & x260 ;
  assign n2437 = ~n2435 & ~n2436 ;
  assign n2438 = ~n2434 & ~n2437 ;
  assign n2439 = n2434 & n2437 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = ~x38 & ~x262 ;
  assign n2442 = x38 & x262 ;
  assign n2443 = ~n2441 & ~n2442 ;
  assign n2444 = ~n2440 & ~n2443 ;
  assign n2445 = n2440 & n2443 ;
  assign n2446 = ~n2444 & ~n2445 ;
  assign n2447 = n2431 & ~n2446 ;
  assign n2448 = ~n2431 & n2446 ;
  assign n2449 = ~n2447 & ~n2448 ;
  assign n2450 = ~x47 & ~x271 ;
  assign n2451 = x47 & x271 ;
  assign n2452 = ~n2450 & ~n2451 ;
  assign n2453 = ~x46 & ~x270 ;
  assign n2454 = x46 & x270 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2456 = ~n2452 & ~n2455 ;
  assign n2457 = n2452 & n2455 ;
  assign n2458 = ~n2456 & ~n2457 ;
  assign n2459 = ~x48 & ~x272 ;
  assign n2460 = x48 & x272 ;
  assign n2461 = ~n2459 & ~n2460 ;
  assign n2462 = ~n2458 & ~n2461 ;
  assign n2463 = n2458 & n2461 ;
  assign n2464 = ~n2462 & ~n2463 ;
  assign n2465 = ~x42 & ~x266 ;
  assign n2466 = x42 & x266 ;
  assign n2467 = ~n2465 & ~n2466 ;
  assign n2468 = ~n2464 & ~n2467 ;
  assign n2469 = n2464 & n2467 ;
  assign n2470 = ~n2468 & ~n2469 ;
  assign n2471 = ~x44 & ~x268 ;
  assign n2472 = x44 & x268 ;
  assign n2473 = ~n2471 & ~n2472 ;
  assign n2474 = ~x43 & ~x267 ;
  assign n2475 = x43 & x267 ;
  assign n2476 = ~n2474 & ~n2475 ;
  assign n2477 = ~n2473 & ~n2476 ;
  assign n2478 = n2473 & n2476 ;
  assign n2479 = ~n2477 & ~n2478 ;
  assign n2480 = ~x45 & ~x269 ;
  assign n2481 = x45 & x269 ;
  assign n2482 = ~n2480 & ~n2481 ;
  assign n2483 = ~n2479 & ~n2482 ;
  assign n2484 = n2479 & n2482 ;
  assign n2485 = ~n2483 & ~n2484 ;
  assign n2486 = n2470 & ~n2485 ;
  assign n2487 = ~n2470 & n2485 ;
  assign n2488 = ~n2486 & ~n2487 ;
  assign n2489 = ~x34 & ~x258 ;
  assign n2490 = x34 & x258 ;
  assign n2491 = ~n2489 & ~n2490 ;
  assign n2492 = n2488 & ~n2491 ;
  assign n2493 = ~n2488 & n2491 ;
  assign n2494 = ~n2492 & ~n2493 ;
  assign n2495 = n2449 & n2494 ;
  assign n2496 = ~n2449 & ~n2494 ;
  assign n2497 = ~n2495 & ~n2496 ;
  assign n2498 = ~n2406 & n2409 ;
  assign n2499 = ~n2410 & ~n2498 ;
  assign n2500 = n2497 & n2499 ;
  assign n2501 = ~n2410 & ~n2500 ;
  assign n2502 = n2404 & ~n2501 ;
  assign n2503 = ~n2429 & ~n2447 ;
  assign n2504 = ~n2418 & ~n2424 ;
  assign n2505 = ~n2503 & n2504 ;
  assign n2506 = n2503 & ~n2504 ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = ~n2439 & ~n2445 ;
  assign n2509 = n2507 & n2508 ;
  assign n2510 = ~n2507 & ~n2508 ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = ~n2468 & ~n2486 ;
  assign n2513 = ~n2457 & ~n2463 ;
  assign n2514 = ~n2512 & n2513 ;
  assign n2515 = n2512 & ~n2513 ;
  assign n2516 = ~n2514 & ~n2515 ;
  assign n2517 = ~n2478 & ~n2484 ;
  assign n2518 = n2516 & n2517 ;
  assign n2519 = ~n2516 & ~n2517 ;
  assign n2520 = ~n2518 & ~n2519 ;
  assign n2521 = ~n2492 & ~n2495 ;
  assign n2522 = n2520 & ~n2521 ;
  assign n2523 = ~n2520 & n2521 ;
  assign n2524 = ~n2522 & ~n2523 ;
  assign n2525 = n2511 & n2524 ;
  assign n2526 = ~n2511 & ~n2524 ;
  assign n2527 = ~n2525 & ~n2526 ;
  assign n2528 = ~n2404 & n2501 ;
  assign n2529 = ~n2502 & ~n2528 ;
  assign n2530 = n2527 & n2529 ;
  assign n2531 = ~n2502 & ~n2530 ;
  assign n2532 = n2402 & ~n2531 ;
  assign n2533 = ~n2514 & ~n2518 ;
  assign n2534 = ~n2522 & ~n2525 ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2536 = n2533 & n2534 ;
  assign n2537 = ~n2535 & ~n2536 ;
  assign n2538 = ~n2505 & ~n2509 ;
  assign n2539 = n2537 & ~n2538 ;
  assign n2540 = ~n2537 & n2538 ;
  assign n2541 = ~n2539 & ~n2540 ;
  assign n2542 = ~n2402 & n2531 ;
  assign n2543 = ~n2532 & ~n2542 ;
  assign n2544 = n2541 & n2543 ;
  assign n2545 = ~n2532 & ~n2544 ;
  assign n2546 = ~n2400 & ~n2545 ;
  assign n2547 = n2400 & n2545 ;
  assign n2548 = ~n2546 & ~n2547 ;
  assign n2549 = ~n2535 & ~n2539 ;
  assign n2550 = n2548 & ~n2549 ;
  assign n2551 = ~n2546 & ~n2550 ;
  assign n2552 = ~n2548 & n2549 ;
  assign n2553 = ~n2550 & ~n2552 ;
  assign n2554 = ~n2541 & ~n2543 ;
  assign n2555 = ~n2544 & ~n2554 ;
  assign n2556 = ~n2497 & ~n2499 ;
  assign n2557 = ~n2500 & ~n2556 ;
  assign n2558 = ~x32 & ~x256 ;
  assign n2559 = x32 & x256 ;
  assign n2560 = ~n2558 & ~n2559 ;
  assign n2561 = ~n2557 & n2560 ;
  assign n2562 = ~n2527 & ~n2529 ;
  assign n2563 = ~n2530 & ~n2562 ;
  assign n2564 = n2561 & ~n2563 ;
  assign n2565 = ~n2555 & n2564 ;
  assign n2566 = ~n2553 & n2565 ;
  assign n2567 = n2551 & n2566 ;
  assign n2568 = n2284 & n2567 ;
  assign n2569 = ~n571 & n2568 ;
  assign n2570 = n560 & ~n566 ;
  assign n2571 = ~n567 & ~n2570 ;
  assign n2572 = ~n2277 & n2279 ;
  assign n2573 = ~n2280 & ~n2572 ;
  assign n2574 = ~n2000 & n2283 ;
  assign n2575 = n1989 & ~n1995 ;
  assign n2576 = ~n1996 & ~n2575 ;
  assign n2577 = ~n1716 & n1999 ;
  assign n2578 = ~n1125 & ~n1146 ;
  assign n2579 = ~n837 & ~n856 ;
  assign n2580 = ~n2578 & ~n2579 ;
  assign n2581 = ~n1148 & n2580 ;
  assign n2582 = ~n1148 & n1431 ;
  assign n2583 = ~n1415 & ~n1430 ;
  assign n2584 = ~n1431 & ~n2583 ;
  assign n2585 = n2581 & ~n2584 ;
  assign n2586 = n1148 & ~n1431 ;
  assign n2587 = n1421 & ~n1427 ;
  assign n2588 = ~n1428 & ~n2587 ;
  assign n2589 = ~n1135 & ~n1139 ;
  assign n2590 = ~n1140 & ~n2589 ;
  assign n2591 = n857 & ~n1147 ;
  assign n2592 = ~n857 & ~n2579 ;
  assign n2593 = ~n1147 & ~n2578 ;
  assign n2594 = n2592 & ~n2593 ;
  assign n2595 = n1127 & ~n1145 ;
  assign n2596 = ~n1146 & ~n2595 ;
  assign n2597 = ~n1140 & ~n1144 ;
  assign n2598 = ~n1145 & ~n2597 ;
  assign n2599 = ~n841 & ~n844 ;
  assign n2600 = ~n845 & ~n2599 ;
  assign n2601 = ~n1130 & n1134 ;
  assign n2602 = ~n1135 & ~n2601 ;
  assign n2603 = ~n2600 & n2602 ;
  assign n2604 = n1139 & n2603 ;
  assign n2605 = ~n845 & ~n849 ;
  assign n2606 = ~n850 & ~n2605 ;
  assign n2607 = ~n2590 & ~n2603 ;
  assign n2608 = ~n2606 & ~n2607 ;
  assign n2609 = ~n2604 & ~n2608 ;
  assign n2610 = n2598 & ~n2609 ;
  assign n2611 = ~n2598 & n2609 ;
  assign n2612 = ~n850 & ~n854 ;
  assign n2613 = ~n855 & ~n2612 ;
  assign n2614 = ~n2611 & ~n2613 ;
  assign n2615 = ~n2610 & ~n2614 ;
  assign n2616 = ~n2596 & n2615 ;
  assign n2617 = n839 & ~n855 ;
  assign n2618 = ~n856 & ~n2617 ;
  assign n2619 = n2596 & ~n2615 ;
  assign n2620 = n2618 & ~n2619 ;
  assign n2621 = ~n2616 & ~n2620 ;
  assign n2622 = ~n2594 & n2621 ;
  assign n2623 = ~n857 & n1147 ;
  assign n2624 = ~n2592 & n2593 ;
  assign n2625 = ~n2623 & ~n2624 ;
  assign n2626 = ~n2622 & n2625 ;
  assign n2627 = ~n2591 & ~n2626 ;
  assign n2628 = ~n2590 & ~n2627 ;
  assign n2629 = ~n2606 & n2627 ;
  assign n2630 = ~n2628 & ~n2629 ;
  assign n2631 = ~n2588 & n2630 ;
  assign n2632 = n1423 & ~n1426 ;
  assign n2633 = ~n1427 & ~n2632 ;
  assign n2634 = ~n2602 & ~n2627 ;
  assign n2635 = ~n2600 & n2627 ;
  assign n2636 = ~n2634 & ~n2635 ;
  assign n2637 = n2633 & ~n2636 ;
  assign n2638 = ~n2631 & n2637 ;
  assign n2639 = n1419 & ~n1428 ;
  assign n2640 = ~n1429 & ~n2639 ;
  assign n2641 = ~n2598 & ~n2627 ;
  assign n2642 = ~n2613 & n2627 ;
  assign n2643 = ~n2641 & ~n2642 ;
  assign n2644 = n2640 & ~n2643 ;
  assign n2645 = n2588 & ~n2630 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = ~n2638 & n2646 ;
  assign n2648 = n1417 & ~n1429 ;
  assign n2649 = ~n1430 & ~n2648 ;
  assign n2650 = ~n2596 & ~n2627 ;
  assign n2651 = ~n2618 & n2627 ;
  assign n2652 = ~n2650 & ~n2651 ;
  assign n2653 = ~n2649 & n2652 ;
  assign n2654 = ~n2640 & n2643 ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = ~n2647 & n2655 ;
  assign n2657 = n2649 & ~n2652 ;
  assign n2658 = ~n2581 & n2584 ;
  assign n2659 = ~n2657 & ~n2658 ;
  assign n2660 = ~n2656 & n2659 ;
  assign n2661 = ~n2586 & ~n2660 ;
  assign n2662 = ~n2585 & n2661 ;
  assign n2663 = ~n2582 & ~n2662 ;
  assign n2664 = n2581 & ~n2663 ;
  assign n2665 = n2584 & ~n2661 ;
  assign n2666 = ~n2664 & ~n2665 ;
  assign n2667 = ~n1432 & n1715 ;
  assign n2668 = n1705 & ~n1711 ;
  assign n2669 = ~n1712 & ~n2668 ;
  assign n2670 = ~n2588 & n2663 ;
  assign n2671 = ~n2630 & ~n2663 ;
  assign n2672 = ~n2670 & ~n2671 ;
  assign n2673 = ~n2669 & n2672 ;
  assign n2674 = n1707 & ~n1710 ;
  assign n2675 = ~n1711 & ~n2674 ;
  assign n2676 = n2636 & ~n2663 ;
  assign n2677 = n2633 & n2663 ;
  assign n2678 = ~n2676 & ~n2677 ;
  assign n2679 = n2675 & n2678 ;
  assign n2680 = ~n2673 & n2679 ;
  assign n2681 = n1703 & ~n1712 ;
  assign n2682 = ~n1713 & ~n2681 ;
  assign n2683 = ~n2640 & n2663 ;
  assign n2684 = ~n2643 & ~n2663 ;
  assign n2685 = ~n2683 & ~n2684 ;
  assign n2686 = n2682 & ~n2685 ;
  assign n2687 = n2669 & ~n2672 ;
  assign n2688 = ~n2686 & ~n2687 ;
  assign n2689 = ~n2680 & n2688 ;
  assign n2690 = n1701 & ~n1713 ;
  assign n2691 = ~n1714 & ~n2690 ;
  assign n2692 = ~n2649 & n2663 ;
  assign n2693 = ~n2652 & ~n2663 ;
  assign n2694 = ~n2692 & ~n2693 ;
  assign n2695 = ~n2691 & n2694 ;
  assign n2696 = ~n2682 & n2685 ;
  assign n2697 = ~n2695 & ~n2696 ;
  assign n2698 = ~n2689 & n2697 ;
  assign n2699 = ~n1699 & ~n1714 ;
  assign n2700 = ~n1715 & ~n2699 ;
  assign n2701 = n2666 & n2700 ;
  assign n2702 = n2691 & ~n2694 ;
  assign n2703 = ~n2701 & ~n2702 ;
  assign n2704 = ~n2698 & n2703 ;
  assign n2705 = n1432 & ~n1715 ;
  assign n2706 = ~n2666 & ~n2700 ;
  assign n2707 = ~n2705 & ~n2706 ;
  assign n2708 = ~n2704 & n2707 ;
  assign n2709 = ~n2667 & ~n2708 ;
  assign n2710 = ~n2666 & ~n2709 ;
  assign n2711 = n2700 & ~n2708 ;
  assign n2712 = ~n2710 & ~n2711 ;
  assign n2713 = ~n1983 & ~n1998 ;
  assign n2714 = ~n1999 & ~n2713 ;
  assign n2715 = ~n2712 & ~n2714 ;
  assign n2716 = n1716 & ~n1999 ;
  assign n2717 = ~n2669 & n2709 ;
  assign n2718 = ~n2672 & ~n2709 ;
  assign n2719 = ~n2717 & ~n2718 ;
  assign n2720 = ~n2576 & n2719 ;
  assign n2721 = n1991 & ~n1994 ;
  assign n2722 = ~n1995 & ~n2721 ;
  assign n2723 = n2678 & ~n2709 ;
  assign n2724 = ~n2675 & n2709 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = n2722 & ~n2725 ;
  assign n2727 = ~n2720 & n2726 ;
  assign n2728 = n1987 & ~n1996 ;
  assign n2729 = ~n1997 & ~n2728 ;
  assign n2730 = n2685 & ~n2709 ;
  assign n2731 = n2682 & n2709 ;
  assign n2732 = ~n2730 & ~n2731 ;
  assign n2733 = n2729 & n2732 ;
  assign n2734 = n2576 & ~n2719 ;
  assign n2735 = ~n2733 & ~n2734 ;
  assign n2736 = ~n2727 & n2735 ;
  assign n2737 = n1985 & ~n1997 ;
  assign n2738 = ~n1998 & ~n2737 ;
  assign n2739 = ~n2691 & n2709 ;
  assign n2740 = ~n2694 & ~n2709 ;
  assign n2741 = ~n2739 & ~n2740 ;
  assign n2742 = ~n2738 & n2741 ;
  assign n2743 = ~n2729 & ~n2732 ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = ~n2736 & n2744 ;
  assign n2746 = n2738 & ~n2741 ;
  assign n2747 = n2712 & n2714 ;
  assign n2748 = ~n2746 & ~n2747 ;
  assign n2749 = ~n2745 & n2748 ;
  assign n2750 = ~n2716 & ~n2749 ;
  assign n2751 = ~n2715 & n2750 ;
  assign n2752 = ~n2577 & ~n2751 ;
  assign n2753 = ~n2576 & n2752 ;
  assign n2754 = ~n2719 & ~n2752 ;
  assign n2755 = ~n2753 & ~n2754 ;
  assign n2756 = ~n2573 & n2755 ;
  assign n2757 = n2273 & ~n2276 ;
  assign n2758 = ~n2277 & ~n2757 ;
  assign n2759 = n2725 & ~n2752 ;
  assign n2760 = n2722 & n2752 ;
  assign n2761 = ~n2759 & ~n2760 ;
  assign n2762 = n2758 & n2761 ;
  assign n2763 = ~n2756 & n2762 ;
  assign n2764 = n2271 & ~n2280 ;
  assign n2765 = ~n2281 & ~n2764 ;
  assign n2766 = ~n2729 & n2752 ;
  assign n2767 = n2732 & ~n2752 ;
  assign n2768 = ~n2766 & ~n2767 ;
  assign n2769 = n2765 & ~n2768 ;
  assign n2770 = n2573 & ~n2755 ;
  assign n2771 = ~n2769 & ~n2770 ;
  assign n2772 = ~n2763 & n2771 ;
  assign n2773 = n2269 & ~n2281 ;
  assign n2774 = ~n2282 & ~n2773 ;
  assign n2775 = ~n2738 & n2752 ;
  assign n2776 = ~n2741 & ~n2752 ;
  assign n2777 = ~n2775 & ~n2776 ;
  assign n2778 = ~n2774 & n2777 ;
  assign n2779 = ~n2765 & n2768 ;
  assign n2780 = ~n2778 & ~n2779 ;
  assign n2781 = ~n2772 & n2780 ;
  assign n2782 = ~n2712 & ~n2752 ;
  assign n2783 = n2714 & ~n2750 ;
  assign n2784 = ~n2782 & ~n2783 ;
  assign n2785 = ~n2267 & ~n2282 ;
  assign n2786 = ~n2283 & ~n2785 ;
  assign n2787 = n2784 & n2786 ;
  assign n2788 = n2774 & ~n2777 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = ~n2781 & n2789 ;
  assign n2791 = n2000 & ~n2283 ;
  assign n2792 = ~n2784 & ~n2786 ;
  assign n2793 = ~n2791 & ~n2792 ;
  assign n2794 = ~n2790 & n2793 ;
  assign n2795 = ~n2574 & ~n2794 ;
  assign n2796 = ~n2573 & n2795 ;
  assign n2797 = ~n2755 & ~n2795 ;
  assign n2798 = ~n2796 & ~n2797 ;
  assign n2799 = ~n2284 & n2567 ;
  assign n2800 = ~n2784 & ~n2795 ;
  assign n2801 = n2786 & ~n2794 ;
  assign n2802 = ~n2800 & ~n2801 ;
  assign n2803 = ~n2551 & ~n2566 ;
  assign n2804 = ~n2567 & ~n2803 ;
  assign n2805 = ~n2802 & ~n2804 ;
  assign n2806 = n2284 & ~n2567 ;
  assign n2807 = ~n2561 & n2563 ;
  assign n2808 = ~n2564 & ~n2807 ;
  assign n2809 = n2798 & ~n2808 ;
  assign n2810 = n2557 & ~n2560 ;
  assign n2811 = ~n2561 & ~n2810 ;
  assign n2812 = n2761 & ~n2795 ;
  assign n2813 = ~n2758 & n2795 ;
  assign n2814 = ~n2812 & ~n2813 ;
  assign n2815 = n2811 & ~n2814 ;
  assign n2816 = ~n2809 & n2815 ;
  assign n2817 = n2555 & ~n2564 ;
  assign n2818 = ~n2565 & ~n2817 ;
  assign n2819 = n2768 & ~n2795 ;
  assign n2820 = n2765 & n2795 ;
  assign n2821 = ~n2819 & ~n2820 ;
  assign n2822 = n2818 & n2821 ;
  assign n2823 = ~n2798 & n2808 ;
  assign n2824 = ~n2822 & ~n2823 ;
  assign n2825 = ~n2816 & n2824 ;
  assign n2826 = n2553 & ~n2565 ;
  assign n2827 = ~n2566 & ~n2826 ;
  assign n2828 = ~n2774 & n2795 ;
  assign n2829 = ~n2777 & ~n2795 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = ~n2827 & n2830 ;
  assign n2832 = ~n2818 & ~n2821 ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2834 = ~n2825 & n2833 ;
  assign n2835 = n2827 & ~n2830 ;
  assign n2836 = n2802 & n2804 ;
  assign n2837 = ~n2835 & ~n2836 ;
  assign n2838 = ~n2834 & n2837 ;
  assign n2839 = ~n2806 & ~n2838 ;
  assign n2840 = ~n2805 & n2839 ;
  assign n2841 = ~n2799 & ~n2840 ;
  assign n2842 = n2798 & ~n2841 ;
  assign n2843 = n2808 & n2841 ;
  assign n2844 = ~n2842 & ~n2843 ;
  assign n2845 = n2571 & n2844 ;
  assign n2846 = n2814 & ~n2841 ;
  assign n2847 = n2811 & n2841 ;
  assign n2848 = n562 & ~n565 ;
  assign n2849 = ~n566 & ~n2848 ;
  assign n2850 = ~n2847 & n2849 ;
  assign n2851 = ~n2846 & n2850 ;
  assign n2852 = ~n2845 & ~n2851 ;
  assign n2853 = ~n2571 & ~n2844 ;
  assign n2854 = n558 & ~n567 ;
  assign n2855 = ~n568 & ~n2854 ;
  assign n2856 = ~n2821 & ~n2841 ;
  assign n2857 = n2818 & n2841 ;
  assign n2858 = ~n2856 & ~n2857 ;
  assign n2859 = ~n2855 & ~n2858 ;
  assign n2860 = ~n2853 & ~n2859 ;
  assign n2861 = ~n2852 & n2860 ;
  assign n2862 = n556 & ~n568 ;
  assign n2863 = ~n569 & ~n2862 ;
  assign n2864 = ~n2827 & n2841 ;
  assign n2865 = ~n2830 & ~n2841 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = n2863 & ~n2866 ;
  assign n2868 = n2855 & n2858 ;
  assign n2869 = ~n2867 & ~n2868 ;
  assign n2870 = ~n2861 & n2869 ;
  assign n2871 = ~n2863 & n2866 ;
  assign n2872 = ~n569 & ~n570 ;
  assign n2873 = ~n571 & ~n2872 ;
  assign n2874 = ~n2802 & ~n2841 ;
  assign n2875 = n2804 & ~n2839 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = ~n2873 & ~n2876 ;
  assign n2878 = ~n2871 & ~n2877 ;
  assign n2879 = ~n2870 & n2878 ;
  assign n2880 = n571 & ~n2568 ;
  assign n2881 = n2873 & n2876 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = ~n2879 & n2882 ;
  assign n2884 = ~n2569 & ~n2883 ;
  assign n2885 = ~x0 & ~n2884 ;
  assign n2886 = ~x32 & n2841 ;
  assign n2887 = ~x192 & ~n2627 ;
  assign n2888 = ~x224 & n2627 ;
  assign n2889 = ~n2887 & ~n2888 ;
  assign n2890 = ~n2663 & ~n2889 ;
  assign n2891 = ~x160 & n2663 ;
  assign n2892 = ~n2890 & ~n2891 ;
  assign n2893 = ~n2709 & n2892 ;
  assign n2894 = x128 & n2709 ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = ~n2752 & ~n2895 ;
  assign n2897 = x96 & n2752 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = ~n2795 & ~n2898 ;
  assign n2900 = x64 & n2795 ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = ~n2841 & n2901 ;
  assign n2903 = ~n2886 & ~n2902 ;
  assign n2904 = n2884 & ~n2903 ;
  assign n2905 = ~n2885 & ~n2904 ;
  assign n2906 = ~x1 & ~n2884 ;
  assign n2907 = ~x33 & n2841 ;
  assign n2908 = ~x193 & ~n2627 ;
  assign n2909 = ~x225 & n2627 ;
  assign n2910 = ~n2908 & ~n2909 ;
  assign n2911 = ~n2663 & ~n2910 ;
  assign n2912 = ~x161 & n2663 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2914 = ~n2709 & n2913 ;
  assign n2915 = x129 & n2709 ;
  assign n2916 = ~n2914 & ~n2915 ;
  assign n2917 = ~n2752 & ~n2916 ;
  assign n2918 = x97 & n2752 ;
  assign n2919 = ~n2917 & ~n2918 ;
  assign n2920 = ~n2795 & ~n2919 ;
  assign n2921 = x65 & n2795 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~n2841 & n2922 ;
  assign n2924 = ~n2907 & ~n2923 ;
  assign n2925 = n2884 & ~n2924 ;
  assign n2926 = ~n2906 & ~n2925 ;
  assign n2927 = ~x2 & ~n2884 ;
  assign n2928 = ~x34 & n2841 ;
  assign n2929 = ~x194 & ~n2627 ;
  assign n2930 = ~x226 & n2627 ;
  assign n2931 = ~n2929 & ~n2930 ;
  assign n2932 = ~n2663 & ~n2931 ;
  assign n2933 = ~x162 & n2663 ;
  assign n2934 = ~n2932 & ~n2933 ;
  assign n2935 = ~n2709 & n2934 ;
  assign n2936 = x130 & n2709 ;
  assign n2937 = ~n2935 & ~n2936 ;
  assign n2938 = ~n2752 & ~n2937 ;
  assign n2939 = x98 & n2752 ;
  assign n2940 = ~n2938 & ~n2939 ;
  assign n2941 = ~n2795 & ~n2940 ;
  assign n2942 = x66 & n2795 ;
  assign n2943 = ~n2941 & ~n2942 ;
  assign n2944 = ~n2841 & n2943 ;
  assign n2945 = ~n2928 & ~n2944 ;
  assign n2946 = n2884 & ~n2945 ;
  assign n2947 = ~n2927 & ~n2946 ;
  assign n2948 = ~x3 & ~n2884 ;
  assign n2949 = ~x35 & n2841 ;
  assign n2950 = ~x195 & ~n2627 ;
  assign n2951 = ~x227 & n2627 ;
  assign n2952 = ~n2950 & ~n2951 ;
  assign n2953 = ~n2663 & ~n2952 ;
  assign n2954 = ~x163 & n2663 ;
  assign n2955 = ~n2953 & ~n2954 ;
  assign n2956 = ~n2709 & n2955 ;
  assign n2957 = x131 & n2709 ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = ~n2752 & ~n2958 ;
  assign n2960 = x99 & n2752 ;
  assign n2961 = ~n2959 & ~n2960 ;
  assign n2962 = ~n2795 & ~n2961 ;
  assign n2963 = x67 & n2795 ;
  assign n2964 = ~n2962 & ~n2963 ;
  assign n2965 = ~n2841 & n2964 ;
  assign n2966 = ~n2949 & ~n2965 ;
  assign n2967 = n2884 & ~n2966 ;
  assign n2968 = ~n2948 & ~n2967 ;
  assign n2969 = ~x4 & ~n2884 ;
  assign n2970 = ~x36 & n2841 ;
  assign n2971 = ~x196 & ~n2627 ;
  assign n2972 = ~x228 & n2627 ;
  assign n2973 = ~n2971 & ~n2972 ;
  assign n2974 = ~n2663 & ~n2973 ;
  assign n2975 = ~x164 & n2663 ;
  assign n2976 = ~n2974 & ~n2975 ;
  assign n2977 = ~n2709 & n2976 ;
  assign n2978 = x132 & n2709 ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = ~n2752 & ~n2979 ;
  assign n2981 = x100 & n2752 ;
  assign n2982 = ~n2980 & ~n2981 ;
  assign n2983 = ~n2795 & ~n2982 ;
  assign n2984 = x68 & n2795 ;
  assign n2985 = ~n2983 & ~n2984 ;
  assign n2986 = ~n2841 & n2985 ;
  assign n2987 = ~n2970 & ~n2986 ;
  assign n2988 = n2884 & ~n2987 ;
  assign n2989 = ~n2969 & ~n2988 ;
  assign n2990 = ~x5 & ~n2884 ;
  assign n2991 = ~x37 & n2841 ;
  assign n2992 = ~x197 & ~n2627 ;
  assign n2993 = ~x229 & n2627 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n2995 = ~n2663 & ~n2994 ;
  assign n2996 = ~x165 & n2663 ;
  assign n2997 = ~n2995 & ~n2996 ;
  assign n2998 = ~n2709 & n2997 ;
  assign n2999 = x133 & n2709 ;
  assign n3000 = ~n2998 & ~n2999 ;
  assign n3001 = ~n2752 & ~n3000 ;
  assign n3002 = x101 & n2752 ;
  assign n3003 = ~n3001 & ~n3002 ;
  assign n3004 = ~n2795 & ~n3003 ;
  assign n3005 = x69 & n2795 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = ~n2841 & n3006 ;
  assign n3008 = ~n2991 & ~n3007 ;
  assign n3009 = n2884 & ~n3008 ;
  assign n3010 = ~n2990 & ~n3009 ;
  assign n3011 = ~x6 & ~n2884 ;
  assign n3012 = ~x38 & n2841 ;
  assign n3013 = ~x198 & ~n2627 ;
  assign n3014 = ~x230 & n2627 ;
  assign n3015 = ~n3013 & ~n3014 ;
  assign n3016 = ~n2663 & ~n3015 ;
  assign n3017 = ~x166 & n2663 ;
  assign n3018 = ~n3016 & ~n3017 ;
  assign n3019 = ~n2709 & n3018 ;
  assign n3020 = x134 & n2709 ;
  assign n3021 = ~n3019 & ~n3020 ;
  assign n3022 = ~n2752 & ~n3021 ;
  assign n3023 = x102 & n2752 ;
  assign n3024 = ~n3022 & ~n3023 ;
  assign n3025 = ~n2795 & ~n3024 ;
  assign n3026 = x70 & n2795 ;
  assign n3027 = ~n3025 & ~n3026 ;
  assign n3028 = ~n2841 & n3027 ;
  assign n3029 = ~n3012 & ~n3028 ;
  assign n3030 = n2884 & ~n3029 ;
  assign n3031 = ~n3011 & ~n3030 ;
  assign n3032 = ~x7 & ~n2884 ;
  assign n3033 = ~x39 & n2841 ;
  assign n3034 = ~x199 & ~n2627 ;
  assign n3035 = ~x231 & n2627 ;
  assign n3036 = ~n3034 & ~n3035 ;
  assign n3037 = ~n2663 & ~n3036 ;
  assign n3038 = ~x167 & n2663 ;
  assign n3039 = ~n3037 & ~n3038 ;
  assign n3040 = ~n2709 & n3039 ;
  assign n3041 = x135 & n2709 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = ~n2752 & ~n3042 ;
  assign n3044 = x103 & n2752 ;
  assign n3045 = ~n3043 & ~n3044 ;
  assign n3046 = ~n2795 & ~n3045 ;
  assign n3047 = x71 & n2795 ;
  assign n3048 = ~n3046 & ~n3047 ;
  assign n3049 = ~n2841 & n3048 ;
  assign n3050 = ~n3033 & ~n3049 ;
  assign n3051 = n2884 & ~n3050 ;
  assign n3052 = ~n3032 & ~n3051 ;
  assign n3053 = ~x8 & ~n2884 ;
  assign n3054 = ~x40 & n2841 ;
  assign n3055 = ~x200 & ~n2627 ;
  assign n3056 = ~x232 & n2627 ;
  assign n3057 = ~n3055 & ~n3056 ;
  assign n3058 = ~n2663 & ~n3057 ;
  assign n3059 = ~x168 & n2663 ;
  assign n3060 = ~n3058 & ~n3059 ;
  assign n3061 = ~n2709 & n3060 ;
  assign n3062 = x136 & n2709 ;
  assign n3063 = ~n3061 & ~n3062 ;
  assign n3064 = ~n2752 & ~n3063 ;
  assign n3065 = x104 & n2752 ;
  assign n3066 = ~n3064 & ~n3065 ;
  assign n3067 = ~n2795 & ~n3066 ;
  assign n3068 = x72 & n2795 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = ~n2841 & n3069 ;
  assign n3071 = ~n3054 & ~n3070 ;
  assign n3072 = n2884 & ~n3071 ;
  assign n3073 = ~n3053 & ~n3072 ;
  assign n3074 = ~x9 & ~n2884 ;
  assign n3075 = ~x41 & n2841 ;
  assign n3076 = ~x201 & ~n2627 ;
  assign n3077 = ~x233 & n2627 ;
  assign n3078 = ~n3076 & ~n3077 ;
  assign n3079 = ~n2663 & ~n3078 ;
  assign n3080 = ~x169 & n2663 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3082 = ~n2709 & n3081 ;
  assign n3083 = x137 & n2709 ;
  assign n3084 = ~n3082 & ~n3083 ;
  assign n3085 = ~n2752 & ~n3084 ;
  assign n3086 = x105 & n2752 ;
  assign n3087 = ~n3085 & ~n3086 ;
  assign n3088 = ~n2795 & ~n3087 ;
  assign n3089 = x73 & n2795 ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = ~n2841 & n3090 ;
  assign n3092 = ~n3075 & ~n3091 ;
  assign n3093 = n2884 & ~n3092 ;
  assign n3094 = ~n3074 & ~n3093 ;
  assign n3095 = ~x10 & ~n2884 ;
  assign n3096 = ~x42 & n2841 ;
  assign n3097 = ~x202 & ~n2627 ;
  assign n3098 = ~x234 & n2627 ;
  assign n3099 = ~n3097 & ~n3098 ;
  assign n3100 = ~n2663 & ~n3099 ;
  assign n3101 = ~x170 & n2663 ;
  assign n3102 = ~n3100 & ~n3101 ;
  assign n3103 = ~n2709 & n3102 ;
  assign n3104 = x138 & n2709 ;
  assign n3105 = ~n3103 & ~n3104 ;
  assign n3106 = ~n2752 & ~n3105 ;
  assign n3107 = x106 & n2752 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = ~n2795 & ~n3108 ;
  assign n3110 = x74 & n2795 ;
  assign n3111 = ~n3109 & ~n3110 ;
  assign n3112 = ~n2841 & n3111 ;
  assign n3113 = ~n3096 & ~n3112 ;
  assign n3114 = n2884 & ~n3113 ;
  assign n3115 = ~n3095 & ~n3114 ;
  assign n3116 = ~x11 & ~n2884 ;
  assign n3117 = ~x43 & n2841 ;
  assign n3118 = ~x203 & ~n2627 ;
  assign n3119 = ~x235 & n2627 ;
  assign n3120 = ~n3118 & ~n3119 ;
  assign n3121 = ~n2663 & ~n3120 ;
  assign n3122 = ~x171 & n2663 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = ~n2709 & n3123 ;
  assign n3125 = x139 & n2709 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = ~n2752 & ~n3126 ;
  assign n3128 = x107 & n2752 ;
  assign n3129 = ~n3127 & ~n3128 ;
  assign n3130 = ~n2795 & ~n3129 ;
  assign n3131 = x75 & n2795 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = ~n2841 & n3132 ;
  assign n3134 = ~n3117 & ~n3133 ;
  assign n3135 = n2884 & ~n3134 ;
  assign n3136 = ~n3116 & ~n3135 ;
  assign n3137 = ~x12 & ~n2884 ;
  assign n3138 = ~x44 & n2841 ;
  assign n3139 = ~x204 & ~n2627 ;
  assign n3140 = ~x236 & n2627 ;
  assign n3141 = ~n3139 & ~n3140 ;
  assign n3142 = ~n2663 & ~n3141 ;
  assign n3143 = ~x172 & n2663 ;
  assign n3144 = ~n3142 & ~n3143 ;
  assign n3145 = ~n2709 & n3144 ;
  assign n3146 = x140 & n2709 ;
  assign n3147 = ~n3145 & ~n3146 ;
  assign n3148 = ~n2752 & ~n3147 ;
  assign n3149 = x108 & n2752 ;
  assign n3150 = ~n3148 & ~n3149 ;
  assign n3151 = ~n2795 & ~n3150 ;
  assign n3152 = x76 & n2795 ;
  assign n3153 = ~n3151 & ~n3152 ;
  assign n3154 = ~n2841 & n3153 ;
  assign n3155 = ~n3138 & ~n3154 ;
  assign n3156 = n2884 & ~n3155 ;
  assign n3157 = ~n3137 & ~n3156 ;
  assign n3158 = ~x13 & ~n2884 ;
  assign n3159 = ~x45 & n2841 ;
  assign n3160 = ~x205 & ~n2627 ;
  assign n3161 = ~x237 & n2627 ;
  assign n3162 = ~n3160 & ~n3161 ;
  assign n3163 = ~n2663 & ~n3162 ;
  assign n3164 = ~x173 & n2663 ;
  assign n3165 = ~n3163 & ~n3164 ;
  assign n3166 = ~n2709 & n3165 ;
  assign n3167 = x141 & n2709 ;
  assign n3168 = ~n3166 & ~n3167 ;
  assign n3169 = ~n2752 & ~n3168 ;
  assign n3170 = x109 & n2752 ;
  assign n3171 = ~n3169 & ~n3170 ;
  assign n3172 = ~n2795 & ~n3171 ;
  assign n3173 = x77 & n2795 ;
  assign n3174 = ~n3172 & ~n3173 ;
  assign n3175 = ~n2841 & n3174 ;
  assign n3176 = ~n3159 & ~n3175 ;
  assign n3177 = n2884 & ~n3176 ;
  assign n3178 = ~n3158 & ~n3177 ;
  assign n3179 = ~x14 & ~n2884 ;
  assign n3180 = ~x46 & n2841 ;
  assign n3181 = ~x206 & ~n2627 ;
  assign n3182 = ~x238 & n2627 ;
  assign n3183 = ~n3181 & ~n3182 ;
  assign n3184 = ~n2663 & ~n3183 ;
  assign n3185 = ~x174 & n2663 ;
  assign n3186 = ~n3184 & ~n3185 ;
  assign n3187 = ~n2709 & n3186 ;
  assign n3188 = x142 & n2709 ;
  assign n3189 = ~n3187 & ~n3188 ;
  assign n3190 = ~n2752 & ~n3189 ;
  assign n3191 = x110 & n2752 ;
  assign n3192 = ~n3190 & ~n3191 ;
  assign n3193 = ~n2795 & ~n3192 ;
  assign n3194 = x78 & n2795 ;
  assign n3195 = ~n3193 & ~n3194 ;
  assign n3196 = ~n2841 & n3195 ;
  assign n3197 = ~n3180 & ~n3196 ;
  assign n3198 = n2884 & ~n3197 ;
  assign n3199 = ~n3179 & ~n3198 ;
  assign n3200 = ~x15 & ~n2884 ;
  assign n3201 = ~x47 & n2841 ;
  assign n3202 = ~x207 & ~n2627 ;
  assign n3203 = ~x239 & n2627 ;
  assign n3204 = ~n3202 & ~n3203 ;
  assign n3205 = ~n2663 & ~n3204 ;
  assign n3206 = ~x175 & n2663 ;
  assign n3207 = ~n3205 & ~n3206 ;
  assign n3208 = ~n2709 & n3207 ;
  assign n3209 = x143 & n2709 ;
  assign n3210 = ~n3208 & ~n3209 ;
  assign n3211 = ~n2752 & ~n3210 ;
  assign n3212 = x111 & n2752 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = ~n2795 & ~n3213 ;
  assign n3215 = x79 & n2795 ;
  assign n3216 = ~n3214 & ~n3215 ;
  assign n3217 = ~n2841 & n3216 ;
  assign n3218 = ~n3201 & ~n3217 ;
  assign n3219 = n2884 & ~n3218 ;
  assign n3220 = ~n3200 & ~n3219 ;
  assign n3221 = ~x16 & ~n2884 ;
  assign n3222 = ~x48 & n2841 ;
  assign n3223 = ~x208 & ~n2627 ;
  assign n3224 = ~x240 & n2627 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = ~n2663 & ~n3225 ;
  assign n3227 = ~x176 & n2663 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = ~n2709 & n3228 ;
  assign n3230 = x144 & n2709 ;
  assign n3231 = ~n3229 & ~n3230 ;
  assign n3232 = ~n2752 & ~n3231 ;
  assign n3233 = x112 & n2752 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3235 = ~n2795 & ~n3234 ;
  assign n3236 = x80 & n2795 ;
  assign n3237 = ~n3235 & ~n3236 ;
  assign n3238 = ~n2841 & n3237 ;
  assign n3239 = ~n3222 & ~n3238 ;
  assign n3240 = n2884 & ~n3239 ;
  assign n3241 = ~n3221 & ~n3240 ;
  assign n3242 = ~x17 & ~n2884 ;
  assign n3243 = ~x49 & n2841 ;
  assign n3244 = ~x209 & ~n2627 ;
  assign n3245 = ~x241 & n2627 ;
  assign n3246 = ~n3244 & ~n3245 ;
  assign n3247 = ~n2663 & ~n3246 ;
  assign n3248 = ~x177 & n2663 ;
  assign n3249 = ~n3247 & ~n3248 ;
  assign n3250 = ~n2709 & n3249 ;
  assign n3251 = x145 & n2709 ;
  assign n3252 = ~n3250 & ~n3251 ;
  assign n3253 = ~n2752 & ~n3252 ;
  assign n3254 = x113 & n2752 ;
  assign n3255 = ~n3253 & ~n3254 ;
  assign n3256 = ~n2795 & ~n3255 ;
  assign n3257 = x81 & n2795 ;
  assign n3258 = ~n3256 & ~n3257 ;
  assign n3259 = ~n2841 & n3258 ;
  assign n3260 = ~n3243 & ~n3259 ;
  assign n3261 = n2884 & ~n3260 ;
  assign n3262 = ~n3242 & ~n3261 ;
  assign n3263 = ~x18 & ~n2884 ;
  assign n3264 = ~x50 & n2841 ;
  assign n3265 = ~x210 & ~n2627 ;
  assign n3266 = ~x242 & n2627 ;
  assign n3267 = ~n3265 & ~n3266 ;
  assign n3268 = ~n2663 & ~n3267 ;
  assign n3269 = ~x178 & n2663 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = ~n2709 & n3270 ;
  assign n3272 = x146 & n2709 ;
  assign n3273 = ~n3271 & ~n3272 ;
  assign n3274 = ~n2752 & ~n3273 ;
  assign n3275 = x114 & n2752 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign n3277 = ~n2795 & ~n3276 ;
  assign n3278 = x82 & n2795 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = ~n2841 & n3279 ;
  assign n3281 = ~n3264 & ~n3280 ;
  assign n3282 = n2884 & ~n3281 ;
  assign n3283 = ~n3263 & ~n3282 ;
  assign n3284 = ~x19 & ~n2884 ;
  assign n3285 = ~x51 & n2841 ;
  assign n3286 = ~x211 & ~n2627 ;
  assign n3287 = ~x243 & n2627 ;
  assign n3288 = ~n3286 & ~n3287 ;
  assign n3289 = ~n2663 & ~n3288 ;
  assign n3290 = ~x179 & n2663 ;
  assign n3291 = ~n3289 & ~n3290 ;
  assign n3292 = ~n2709 & n3291 ;
  assign n3293 = x147 & n2709 ;
  assign n3294 = ~n3292 & ~n3293 ;
  assign n3295 = ~n2752 & ~n3294 ;
  assign n3296 = x115 & n2752 ;
  assign n3297 = ~n3295 & ~n3296 ;
  assign n3298 = ~n2795 & ~n3297 ;
  assign n3299 = x83 & n2795 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = ~n2841 & n3300 ;
  assign n3302 = ~n3285 & ~n3301 ;
  assign n3303 = n2884 & ~n3302 ;
  assign n3304 = ~n3284 & ~n3303 ;
  assign n3305 = ~x20 & ~n2884 ;
  assign n3306 = ~x52 & n2841 ;
  assign n3307 = ~x212 & ~n2627 ;
  assign n3308 = ~x244 & n2627 ;
  assign n3309 = ~n3307 & ~n3308 ;
  assign n3310 = ~n2663 & ~n3309 ;
  assign n3311 = ~x180 & n2663 ;
  assign n3312 = ~n3310 & ~n3311 ;
  assign n3313 = ~n2709 & n3312 ;
  assign n3314 = x148 & n2709 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3316 = ~n2752 & ~n3315 ;
  assign n3317 = x116 & n2752 ;
  assign n3318 = ~n3316 & ~n3317 ;
  assign n3319 = ~n2795 & ~n3318 ;
  assign n3320 = x84 & n2795 ;
  assign n3321 = ~n3319 & ~n3320 ;
  assign n3322 = ~n2841 & n3321 ;
  assign n3323 = ~n3306 & ~n3322 ;
  assign n3324 = n2884 & ~n3323 ;
  assign n3325 = ~n3305 & ~n3324 ;
  assign n3326 = ~x21 & ~n2884 ;
  assign n3327 = ~x53 & n2841 ;
  assign n3328 = ~x213 & ~n2627 ;
  assign n3329 = ~x245 & n2627 ;
  assign n3330 = ~n3328 & ~n3329 ;
  assign n3331 = ~n2663 & ~n3330 ;
  assign n3332 = ~x181 & n2663 ;
  assign n3333 = ~n3331 & ~n3332 ;
  assign n3334 = ~n2709 & n3333 ;
  assign n3335 = x149 & n2709 ;
  assign n3336 = ~n3334 & ~n3335 ;
  assign n3337 = ~n2752 & ~n3336 ;
  assign n3338 = x117 & n2752 ;
  assign n3339 = ~n3337 & ~n3338 ;
  assign n3340 = ~n2795 & ~n3339 ;
  assign n3341 = x85 & n2795 ;
  assign n3342 = ~n3340 & ~n3341 ;
  assign n3343 = ~n2841 & n3342 ;
  assign n3344 = ~n3327 & ~n3343 ;
  assign n3345 = n2884 & ~n3344 ;
  assign n3346 = ~n3326 & ~n3345 ;
  assign n3347 = ~x22 & ~n2884 ;
  assign n3348 = ~x54 & n2841 ;
  assign n3349 = ~x214 & ~n2627 ;
  assign n3350 = ~x246 & n2627 ;
  assign n3351 = ~n3349 & ~n3350 ;
  assign n3352 = ~n2663 & ~n3351 ;
  assign n3353 = ~x182 & n2663 ;
  assign n3354 = ~n3352 & ~n3353 ;
  assign n3355 = ~n2709 & n3354 ;
  assign n3356 = x150 & n2709 ;
  assign n3357 = ~n3355 & ~n3356 ;
  assign n3358 = ~n2752 & ~n3357 ;
  assign n3359 = x118 & n2752 ;
  assign n3360 = ~n3358 & ~n3359 ;
  assign n3361 = ~n2795 & ~n3360 ;
  assign n3362 = x86 & n2795 ;
  assign n3363 = ~n3361 & ~n3362 ;
  assign n3364 = ~n2841 & n3363 ;
  assign n3365 = ~n3348 & ~n3364 ;
  assign n3366 = n2884 & ~n3365 ;
  assign n3367 = ~n3347 & ~n3366 ;
  assign n3368 = ~x23 & ~n2884 ;
  assign n3369 = ~x55 & n2841 ;
  assign n3370 = ~x215 & ~n2627 ;
  assign n3371 = ~x247 & n2627 ;
  assign n3372 = ~n3370 & ~n3371 ;
  assign n3373 = ~n2663 & ~n3372 ;
  assign n3374 = ~x183 & n2663 ;
  assign n3375 = ~n3373 & ~n3374 ;
  assign n3376 = ~n2709 & n3375 ;
  assign n3377 = x151 & n2709 ;
  assign n3378 = ~n3376 & ~n3377 ;
  assign n3379 = ~n2752 & ~n3378 ;
  assign n3380 = x119 & n2752 ;
  assign n3381 = ~n3379 & ~n3380 ;
  assign n3382 = ~n2795 & ~n3381 ;
  assign n3383 = x87 & n2795 ;
  assign n3384 = ~n3382 & ~n3383 ;
  assign n3385 = ~n2841 & n3384 ;
  assign n3386 = ~n3369 & ~n3385 ;
  assign n3387 = n2884 & ~n3386 ;
  assign n3388 = ~n3368 & ~n3387 ;
  assign n3389 = ~x24 & ~n2884 ;
  assign n3390 = ~x56 & n2841 ;
  assign n3391 = ~x216 & ~n2627 ;
  assign n3392 = ~x248 & n2627 ;
  assign n3393 = ~n3391 & ~n3392 ;
  assign n3394 = ~n2663 & ~n3393 ;
  assign n3395 = ~x184 & n2663 ;
  assign n3396 = ~n3394 & ~n3395 ;
  assign n3397 = ~n2709 & n3396 ;
  assign n3398 = x152 & n2709 ;
  assign n3399 = ~n3397 & ~n3398 ;
  assign n3400 = ~n2752 & ~n3399 ;
  assign n3401 = x120 & n2752 ;
  assign n3402 = ~n3400 & ~n3401 ;
  assign n3403 = ~n2795 & ~n3402 ;
  assign n3404 = x88 & n2795 ;
  assign n3405 = ~n3403 & ~n3404 ;
  assign n3406 = ~n2841 & n3405 ;
  assign n3407 = ~n3390 & ~n3406 ;
  assign n3408 = n2884 & ~n3407 ;
  assign n3409 = ~n3389 & ~n3408 ;
  assign n3410 = ~x25 & ~n2884 ;
  assign n3411 = ~x57 & n2841 ;
  assign n3412 = ~x217 & ~n2627 ;
  assign n3413 = ~x249 & n2627 ;
  assign n3414 = ~n3412 & ~n3413 ;
  assign n3415 = ~n2663 & ~n3414 ;
  assign n3416 = ~x185 & n2663 ;
  assign n3417 = ~n3415 & ~n3416 ;
  assign n3418 = ~n2709 & n3417 ;
  assign n3419 = x153 & n2709 ;
  assign n3420 = ~n3418 & ~n3419 ;
  assign n3421 = ~n2752 & ~n3420 ;
  assign n3422 = x121 & n2752 ;
  assign n3423 = ~n3421 & ~n3422 ;
  assign n3424 = ~n2795 & ~n3423 ;
  assign n3425 = x89 & n2795 ;
  assign n3426 = ~n3424 & ~n3425 ;
  assign n3427 = ~n2841 & n3426 ;
  assign n3428 = ~n3411 & ~n3427 ;
  assign n3429 = n2884 & ~n3428 ;
  assign n3430 = ~n3410 & ~n3429 ;
  assign n3431 = ~x26 & ~n2884 ;
  assign n3432 = ~x58 & n2841 ;
  assign n3433 = ~x218 & ~n2627 ;
  assign n3434 = ~x250 & n2627 ;
  assign n3435 = ~n3433 & ~n3434 ;
  assign n3436 = ~n2663 & ~n3435 ;
  assign n3437 = ~x186 & n2663 ;
  assign n3438 = ~n3436 & ~n3437 ;
  assign n3439 = ~n2709 & n3438 ;
  assign n3440 = x154 & n2709 ;
  assign n3441 = ~n3439 & ~n3440 ;
  assign n3442 = ~n2752 & ~n3441 ;
  assign n3443 = x122 & n2752 ;
  assign n3444 = ~n3442 & ~n3443 ;
  assign n3445 = ~n2795 & ~n3444 ;
  assign n3446 = x90 & n2795 ;
  assign n3447 = ~n3445 & ~n3446 ;
  assign n3448 = ~n2841 & n3447 ;
  assign n3449 = ~n3432 & ~n3448 ;
  assign n3450 = n2884 & ~n3449 ;
  assign n3451 = ~n3431 & ~n3450 ;
  assign n3452 = ~x27 & ~n2884 ;
  assign n3453 = ~x59 & n2841 ;
  assign n3454 = ~x219 & ~n2627 ;
  assign n3455 = ~x251 & n2627 ;
  assign n3456 = ~n3454 & ~n3455 ;
  assign n3457 = ~n2663 & ~n3456 ;
  assign n3458 = ~x187 & n2663 ;
  assign n3459 = ~n3457 & ~n3458 ;
  assign n3460 = ~n2709 & n3459 ;
  assign n3461 = x155 & n2709 ;
  assign n3462 = ~n3460 & ~n3461 ;
  assign n3463 = ~n2752 & ~n3462 ;
  assign n3464 = x123 & n2752 ;
  assign n3465 = ~n3463 & ~n3464 ;
  assign n3466 = ~n2795 & ~n3465 ;
  assign n3467 = x91 & n2795 ;
  assign n3468 = ~n3466 & ~n3467 ;
  assign n3469 = ~n2841 & n3468 ;
  assign n3470 = ~n3453 & ~n3469 ;
  assign n3471 = n2884 & ~n3470 ;
  assign n3472 = ~n3452 & ~n3471 ;
  assign n3473 = ~x28 & ~n2884 ;
  assign n3474 = ~x60 & n2841 ;
  assign n3475 = ~x220 & ~n2627 ;
  assign n3476 = ~x252 & n2627 ;
  assign n3477 = ~n3475 & ~n3476 ;
  assign n3478 = ~n2663 & ~n3477 ;
  assign n3479 = ~x188 & n2663 ;
  assign n3480 = ~n3478 & ~n3479 ;
  assign n3481 = ~n2709 & n3480 ;
  assign n3482 = x156 & n2709 ;
  assign n3483 = ~n3481 & ~n3482 ;
  assign n3484 = ~n2752 & ~n3483 ;
  assign n3485 = x124 & n2752 ;
  assign n3486 = ~n3484 & ~n3485 ;
  assign n3487 = ~n2795 & ~n3486 ;
  assign n3488 = x92 & n2795 ;
  assign n3489 = ~n3487 & ~n3488 ;
  assign n3490 = ~n2841 & n3489 ;
  assign n3491 = ~n3474 & ~n3490 ;
  assign n3492 = n2884 & ~n3491 ;
  assign n3493 = ~n3473 & ~n3492 ;
  assign n3494 = ~x29 & ~n2884 ;
  assign n3495 = ~x61 & n2841 ;
  assign n3496 = ~x221 & ~n2627 ;
  assign n3497 = ~x253 & n2627 ;
  assign n3498 = ~n3496 & ~n3497 ;
  assign n3499 = ~n2663 & ~n3498 ;
  assign n3500 = ~x189 & n2663 ;
  assign n3501 = ~n3499 & ~n3500 ;
  assign n3502 = ~n2709 & n3501 ;
  assign n3503 = x157 & n2709 ;
  assign n3504 = ~n3502 & ~n3503 ;
  assign n3505 = ~n2752 & ~n3504 ;
  assign n3506 = x125 & n2752 ;
  assign n3507 = ~n3505 & ~n3506 ;
  assign n3508 = ~n2795 & ~n3507 ;
  assign n3509 = x93 & n2795 ;
  assign n3510 = ~n3508 & ~n3509 ;
  assign n3511 = ~n2841 & n3510 ;
  assign n3512 = ~n3495 & ~n3511 ;
  assign n3513 = n2884 & ~n3512 ;
  assign n3514 = ~n3494 & ~n3513 ;
  assign n3515 = ~x30 & ~n2884 ;
  assign n3516 = ~x62 & n2841 ;
  assign n3517 = ~x222 & ~n2627 ;
  assign n3518 = ~x254 & n2627 ;
  assign n3519 = ~n3517 & ~n3518 ;
  assign n3520 = ~n2663 & ~n3519 ;
  assign n3521 = ~x190 & n2663 ;
  assign n3522 = ~n3520 & ~n3521 ;
  assign n3523 = ~n2709 & n3522 ;
  assign n3524 = x158 & n2709 ;
  assign n3525 = ~n3523 & ~n3524 ;
  assign n3526 = ~n2752 & ~n3525 ;
  assign n3527 = x126 & n2752 ;
  assign n3528 = ~n3526 & ~n3527 ;
  assign n3529 = ~n2795 & ~n3528 ;
  assign n3530 = x94 & n2795 ;
  assign n3531 = ~n3529 & ~n3530 ;
  assign n3532 = ~n2841 & n3531 ;
  assign n3533 = ~n3516 & ~n3532 ;
  assign n3534 = n2884 & ~n3533 ;
  assign n3535 = ~n3515 & ~n3534 ;
  assign n3536 = ~x31 & ~n2884 ;
  assign n3537 = ~x63 & n2841 ;
  assign n3538 = ~x223 & ~n2627 ;
  assign n3539 = ~x255 & n2627 ;
  assign n3540 = ~n3538 & ~n3539 ;
  assign n3541 = ~n2663 & ~n3540 ;
  assign n3542 = ~x191 & n2663 ;
  assign n3543 = ~n3541 & ~n3542 ;
  assign n3544 = ~n2709 & n3543 ;
  assign n3545 = x159 & n2709 ;
  assign n3546 = ~n3544 & ~n3545 ;
  assign n3547 = ~n2752 & ~n3546 ;
  assign n3548 = x127 & n2752 ;
  assign n3549 = ~n3547 & ~n3548 ;
  assign n3550 = ~n2795 & ~n3549 ;
  assign n3551 = x95 & n2795 ;
  assign n3552 = ~n3550 & ~n3551 ;
  assign n3553 = ~n2841 & n3552 ;
  assign n3554 = ~n3537 & ~n3553 ;
  assign n3555 = n2884 & ~n3554 ;
  assign n3556 = ~n3536 & ~n3555 ;
  assign y0 = n2905 ;
  assign y1 = n2926 ;
  assign y2 = n2947 ;
  assign y3 = n2968 ;
  assign y4 = n2989 ;
  assign y5 = n3010 ;
  assign y6 = n3031 ;
  assign y7 = n3052 ;
  assign y8 = n3073 ;
  assign y9 = n3094 ;
  assign y10 = n3115 ;
  assign y11 = n3136 ;
  assign y12 = n3157 ;
  assign y13 = n3178 ;
  assign y14 = n3199 ;
  assign y15 = n3220 ;
  assign y16 = n3241 ;
  assign y17 = n3262 ;
  assign y18 = n3283 ;
  assign y19 = n3304 ;
  assign y20 = n3325 ;
  assign y21 = n3346 ;
  assign y22 = n3367 ;
  assign y23 = n3388 ;
  assign y24 = n3409 ;
  assign y25 = n3430 ;
  assign y26 = n3451 ;
  assign y27 = n3472 ;
  assign y28 = n3493 ;
  assign y29 = n3514 ;
  assign y30 = n3535 ;
  assign y31 = n3556 ;
endmodule
